//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for sb_2_ -----
module sb_2_(config_enable,
             prog_reset,
             prog_clk,
             chany_top_in,
             top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_,
             top_right_grid_left_width_0_height_0_subtile_4__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_5__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_6__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_7__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_8__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_9__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_10__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_11__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_12__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_13__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_14__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_15__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_16__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_17__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_18__pin_out_0_,
             top_right_grid_left_width_0_height_0_subtile_19__pin_out_0_,
             chanx_right_in,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_,
             right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_,
             chany_bottom_in,
             bottom_right_grid_left_width_0_height_0_subtile_4__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_5__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_6__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_7__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_8__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_9__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_10__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_11__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_12__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_13__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_14__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_15__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_16__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_17__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_18__pin_out_0_,
             bottom_right_grid_left_width_0_height_0_subtile_19__pin_out_0_,
             bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_,
             bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_,
             bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_,
             bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_,
             bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_,
             bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_,
             bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_,
             bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_,
             chanx_left_in,
             ccff_head,
             chany_top_out,
             chanx_right_out,
             chany_bottom_out,
             chanx_left_out,
             ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:63] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_8__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_9__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_10__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_11__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_12__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_13__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_14__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_15__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_16__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_17__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_18__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_19__pin_out_0_;
//----- INPUT PORTS -----
input [0:63] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_;
//----- INPUT PORTS -----
input [0:63] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_8__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_9__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_10__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_11__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_12__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_13__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_14__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_15__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_16__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_17__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_18__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_19__pin_out_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:63] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:63] chany_top_out;
//----- OUTPUT PORTS -----
output [0:63] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:63] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:63] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] clk_mux_size3_0_sram;
wire [0:1] clk_mux_size3_0_sram_inv;
wire [0:1] clk_mux_size3_10_sram;
wire [0:1] clk_mux_size3_10_sram_inv;
wire [0:1] clk_mux_size3_11_sram;
wire [0:1] clk_mux_size3_11_sram_inv;
wire [0:1] clk_mux_size3_12_sram;
wire [0:1] clk_mux_size3_12_sram_inv;
wire [0:1] clk_mux_size3_13_sram;
wire [0:1] clk_mux_size3_13_sram_inv;
wire [0:1] clk_mux_size3_14_sram;
wire [0:1] clk_mux_size3_14_sram_inv;
wire [0:1] clk_mux_size3_15_sram;
wire [0:1] clk_mux_size3_15_sram_inv;
wire [0:1] clk_mux_size3_16_sram;
wire [0:1] clk_mux_size3_16_sram_inv;
wire [0:1] clk_mux_size3_17_sram;
wire [0:1] clk_mux_size3_17_sram_inv;
wire [0:1] clk_mux_size3_18_sram;
wire [0:1] clk_mux_size3_18_sram_inv;
wire [0:1] clk_mux_size3_19_sram;
wire [0:1] clk_mux_size3_19_sram_inv;
wire [0:1] clk_mux_size3_1_sram;
wire [0:1] clk_mux_size3_1_sram_inv;
wire [0:1] clk_mux_size3_20_sram;
wire [0:1] clk_mux_size3_20_sram_inv;
wire [0:1] clk_mux_size3_21_sram;
wire [0:1] clk_mux_size3_21_sram_inv;
wire [0:1] clk_mux_size3_22_sram;
wire [0:1] clk_mux_size3_22_sram_inv;
wire [0:1] clk_mux_size3_23_sram;
wire [0:1] clk_mux_size3_23_sram_inv;
wire [0:1] clk_mux_size3_24_sram;
wire [0:1] clk_mux_size3_24_sram_inv;
wire [0:1] clk_mux_size3_25_sram;
wire [0:1] clk_mux_size3_25_sram_inv;
wire [0:1] clk_mux_size3_26_sram;
wire [0:1] clk_mux_size3_26_sram_inv;
wire [0:1] clk_mux_size3_27_sram;
wire [0:1] clk_mux_size3_27_sram_inv;
wire [0:1] clk_mux_size3_28_sram;
wire [0:1] clk_mux_size3_28_sram_inv;
wire [0:1] clk_mux_size3_29_sram;
wire [0:1] clk_mux_size3_29_sram_inv;
wire [0:1] clk_mux_size3_2_sram;
wire [0:1] clk_mux_size3_2_sram_inv;
wire [0:1] clk_mux_size3_30_sram;
wire [0:1] clk_mux_size3_30_sram_inv;
wire [0:1] clk_mux_size3_31_sram;
wire [0:1] clk_mux_size3_31_sram_inv;
wire [0:1] clk_mux_size3_32_sram;
wire [0:1] clk_mux_size3_32_sram_inv;
wire [0:1] clk_mux_size3_33_sram;
wire [0:1] clk_mux_size3_33_sram_inv;
wire [0:1] clk_mux_size3_34_sram;
wire [0:1] clk_mux_size3_34_sram_inv;
wire [0:1] clk_mux_size3_35_sram;
wire [0:1] clk_mux_size3_35_sram_inv;
wire [0:1] clk_mux_size3_36_sram;
wire [0:1] clk_mux_size3_36_sram_inv;
wire [0:1] clk_mux_size3_37_sram;
wire [0:1] clk_mux_size3_37_sram_inv;
wire [0:1] clk_mux_size3_38_sram;
wire [0:1] clk_mux_size3_38_sram_inv;
wire [0:1] clk_mux_size3_39_sram;
wire [0:1] clk_mux_size3_39_sram_inv;
wire [0:1] clk_mux_size3_3_sram;
wire [0:1] clk_mux_size3_3_sram_inv;
wire [0:1] clk_mux_size3_40_sram;
wire [0:1] clk_mux_size3_40_sram_inv;
wire [0:1] clk_mux_size3_41_sram;
wire [0:1] clk_mux_size3_41_sram_inv;
wire [0:1] clk_mux_size3_42_sram;
wire [0:1] clk_mux_size3_42_sram_inv;
wire [0:1] clk_mux_size3_43_sram;
wire [0:1] clk_mux_size3_43_sram_inv;
wire [0:1] clk_mux_size3_44_sram;
wire [0:1] clk_mux_size3_44_sram_inv;
wire [0:1] clk_mux_size3_45_sram;
wire [0:1] clk_mux_size3_45_sram_inv;
wire [0:1] clk_mux_size3_46_sram;
wire [0:1] clk_mux_size3_46_sram_inv;
wire [0:1] clk_mux_size3_47_sram;
wire [0:1] clk_mux_size3_47_sram_inv;
wire [0:1] clk_mux_size3_48_sram;
wire [0:1] clk_mux_size3_48_sram_inv;
wire [0:1] clk_mux_size3_49_sram;
wire [0:1] clk_mux_size3_49_sram_inv;
wire [0:1] clk_mux_size3_4_sram;
wire [0:1] clk_mux_size3_4_sram_inv;
wire [0:1] clk_mux_size3_50_sram;
wire [0:1] clk_mux_size3_50_sram_inv;
wire [0:1] clk_mux_size3_51_sram;
wire [0:1] clk_mux_size3_51_sram_inv;
wire [0:1] clk_mux_size3_52_sram;
wire [0:1] clk_mux_size3_52_sram_inv;
wire [0:1] clk_mux_size3_53_sram;
wire [0:1] clk_mux_size3_53_sram_inv;
wire [0:1] clk_mux_size3_54_sram;
wire [0:1] clk_mux_size3_54_sram_inv;
wire [0:1] clk_mux_size3_55_sram;
wire [0:1] clk_mux_size3_55_sram_inv;
wire [0:1] clk_mux_size3_56_sram;
wire [0:1] clk_mux_size3_56_sram_inv;
wire [0:1] clk_mux_size3_57_sram;
wire [0:1] clk_mux_size3_57_sram_inv;
wire [0:1] clk_mux_size3_58_sram;
wire [0:1] clk_mux_size3_58_sram_inv;
wire [0:1] clk_mux_size3_59_sram;
wire [0:1] clk_mux_size3_59_sram_inv;
wire [0:1] clk_mux_size3_5_sram;
wire [0:1] clk_mux_size3_5_sram_inv;
wire [0:1] clk_mux_size3_60_sram;
wire [0:1] clk_mux_size3_60_sram_inv;
wire [0:1] clk_mux_size3_61_sram;
wire [0:1] clk_mux_size3_61_sram_inv;
wire [0:1] clk_mux_size3_62_sram;
wire [0:1] clk_mux_size3_62_sram_inv;
wire [0:1] clk_mux_size3_63_sram;
wire [0:1] clk_mux_size3_63_sram_inv;
wire [0:1] clk_mux_size3_64_sram;
wire [0:1] clk_mux_size3_64_sram_inv;
wire [0:1] clk_mux_size3_65_sram;
wire [0:1] clk_mux_size3_65_sram_inv;
wire [0:1] clk_mux_size3_66_sram;
wire [0:1] clk_mux_size3_66_sram_inv;
wire [0:1] clk_mux_size3_67_sram;
wire [0:1] clk_mux_size3_67_sram_inv;
wire [0:1] clk_mux_size3_68_sram;
wire [0:1] clk_mux_size3_68_sram_inv;
wire [0:1] clk_mux_size3_69_sram;
wire [0:1] clk_mux_size3_69_sram_inv;
wire [0:1] clk_mux_size3_6_sram;
wire [0:1] clk_mux_size3_6_sram_inv;
wire [0:1] clk_mux_size3_70_sram;
wire [0:1] clk_mux_size3_70_sram_inv;
wire [0:1] clk_mux_size3_71_sram;
wire [0:1] clk_mux_size3_71_sram_inv;
wire [0:1] clk_mux_size3_72_sram;
wire [0:1] clk_mux_size3_72_sram_inv;
wire [0:1] clk_mux_size3_73_sram;
wire [0:1] clk_mux_size3_73_sram_inv;
wire [0:1] clk_mux_size3_74_sram;
wire [0:1] clk_mux_size3_74_sram_inv;
wire [0:1] clk_mux_size3_75_sram;
wire [0:1] clk_mux_size3_75_sram_inv;
wire [0:1] clk_mux_size3_76_sram;
wire [0:1] clk_mux_size3_76_sram_inv;
wire [0:1] clk_mux_size3_77_sram;
wire [0:1] clk_mux_size3_77_sram_inv;
wire [0:1] clk_mux_size3_78_sram;
wire [0:1] clk_mux_size3_78_sram_inv;
wire [0:1] clk_mux_size3_79_sram;
wire [0:1] clk_mux_size3_79_sram_inv;
wire [0:1] clk_mux_size3_7_sram;
wire [0:1] clk_mux_size3_7_sram_inv;
wire [0:1] clk_mux_size3_80_sram;
wire [0:1] clk_mux_size3_80_sram_inv;
wire [0:1] clk_mux_size3_81_sram;
wire [0:1] clk_mux_size3_81_sram_inv;
wire [0:1] clk_mux_size3_82_sram;
wire [0:1] clk_mux_size3_82_sram_inv;
wire [0:1] clk_mux_size3_83_sram;
wire [0:1] clk_mux_size3_83_sram_inv;
wire [0:1] clk_mux_size3_84_sram;
wire [0:1] clk_mux_size3_84_sram_inv;
wire [0:1] clk_mux_size3_85_sram;
wire [0:1] clk_mux_size3_85_sram_inv;
wire [0:1] clk_mux_size3_86_sram;
wire [0:1] clk_mux_size3_86_sram_inv;
wire [0:1] clk_mux_size3_87_sram;
wire [0:1] clk_mux_size3_87_sram_inv;
wire [0:1] clk_mux_size3_88_sram;
wire [0:1] clk_mux_size3_88_sram_inv;
wire [0:1] clk_mux_size3_89_sram;
wire [0:1] clk_mux_size3_89_sram_inv;
wire [0:1] clk_mux_size3_8_sram;
wire [0:1] clk_mux_size3_8_sram_inv;
wire [0:1] clk_mux_size3_90_sram;
wire [0:1] clk_mux_size3_90_sram_inv;
wire [0:1] clk_mux_size3_91_sram;
wire [0:1] clk_mux_size3_91_sram_inv;
wire [0:1] clk_mux_size3_92_sram;
wire [0:1] clk_mux_size3_92_sram_inv;
wire [0:1] clk_mux_size3_93_sram;
wire [0:1] clk_mux_size3_93_sram_inv;
wire [0:1] clk_mux_size3_94_sram;
wire [0:1] clk_mux_size3_94_sram_inv;
wire [0:1] clk_mux_size3_95_sram;
wire [0:1] clk_mux_size3_95_sram_inv;
wire [0:1] clk_mux_size3_9_sram;
wire [0:1] clk_mux_size3_9_sram_inv;
wire [0:407] sb_2__config_group_mem_size408_0_mem_out;
wire [0:407] sb_2__config_group_mem_size408_0_mem_outb;
wire [0:3] sb_mux_size10_0_sram;
wire [0:3] sb_mux_size10_0_sram_inv;
wire [0:3] sb_mux_size10_1_sram;
wire [0:3] sb_mux_size10_1_sram_inv;
wire [0:3] sb_mux_size10_2_sram;
wire [0:3] sb_mux_size10_2_sram_inv;
wire [0:3] sb_mux_size10_3_sram;
wire [0:3] sb_mux_size10_3_sram_inv;
wire [0:3] sb_mux_size10_4_sram;
wire [0:3] sb_mux_size10_4_sram_inv;
wire [0:3] sb_mux_size10_5_sram;
wire [0:3] sb_mux_size10_5_sram_inv;
wire [0:3] sb_mux_size10_6_sram;
wire [0:3] sb_mux_size10_6_sram_inv;
wire [0:3] sb_mux_size10_7_sram;
wire [0:3] sb_mux_size10_7_sram_inv;
wire [0:3] sb_mux_size11_0_sram;
wire [0:3] sb_mux_size11_0_sram_inv;
wire [0:3] sb_mux_size11_10_sram;
wire [0:3] sb_mux_size11_10_sram_inv;
wire [0:3] sb_mux_size11_11_sram;
wire [0:3] sb_mux_size11_11_sram_inv;
wire [0:3] sb_mux_size11_12_sram;
wire [0:3] sb_mux_size11_12_sram_inv;
wire [0:3] sb_mux_size11_13_sram;
wire [0:3] sb_mux_size11_13_sram_inv;
wire [0:3] sb_mux_size11_1_sram;
wire [0:3] sb_mux_size11_1_sram_inv;
wire [0:3] sb_mux_size11_2_sram;
wire [0:3] sb_mux_size11_2_sram_inv;
wire [0:3] sb_mux_size11_3_sram;
wire [0:3] sb_mux_size11_3_sram_inv;
wire [0:3] sb_mux_size11_4_sram;
wire [0:3] sb_mux_size11_4_sram_inv;
wire [0:3] sb_mux_size11_5_sram;
wire [0:3] sb_mux_size11_5_sram_inv;
wire [0:3] sb_mux_size11_6_sram;
wire [0:3] sb_mux_size11_6_sram_inv;
wire [0:3] sb_mux_size11_7_sram;
wire [0:3] sb_mux_size11_7_sram_inv;
wire [0:3] sb_mux_size11_8_sram;
wire [0:3] sb_mux_size11_8_sram_inv;
wire [0:3] sb_mux_size11_9_sram;
wire [0:3] sb_mux_size11_9_sram_inv;
wire [0:2] sb_mux_size7_0_sram;
wire [0:2] sb_mux_size7_0_sram_inv;
wire [0:2] sb_mux_size7_1_sram;
wire [0:2] sb_mux_size7_1_sram_inv;
wire [0:2] sb_mux_size7_2_sram;
wire [0:2] sb_mux_size7_2_sram_inv;
wire [0:2] sb_mux_size7_3_sram;
wire [0:2] sb_mux_size7_3_sram_inv;
wire [0:2] sb_mux_size7_4_sram;
wire [0:2] sb_mux_size7_4_sram_inv;
wire [0:2] sb_mux_size7_5_sram;
wire [0:2] sb_mux_size7_5_sram_inv;
wire [0:2] sb_mux_size7_6_sram;
wire [0:2] sb_mux_size7_6_sram_inv;
wire [0:2] sb_mux_size7_7_sram;
wire [0:2] sb_mux_size7_7_sram_inv;
wire [0:3] sb_mux_size8_0_sram;
wire [0:3] sb_mux_size8_0_sram_inv;
wire [0:3] sb_mux_size8_1_sram;
wire [0:3] sb_mux_size8_1_sram_inv;
wire [0:3] sb_mux_size8_2_sram;
wire [0:3] sb_mux_size8_2_sram_inv;
wire [0:3] sb_mux_size8_3_sram;
wire [0:3] sb_mux_size8_3_sram_inv;
wire [0:3] sb_mux_size8_4_sram;
wire [0:3] sb_mux_size8_4_sram_inv;
wire [0:3] sb_mux_size8_5_sram;
wire [0:3] sb_mux_size8_5_sram_inv;
wire [0:3] sb_mux_size8_6_sram;
wire [0:3] sb_mux_size8_6_sram_inv;
wire [0:3] sb_mux_size8_7_sram;
wire [0:3] sb_mux_size8_7_sram_inv;
wire [0:3] sb_mux_size9_0_sram;
wire [0:3] sb_mux_size9_0_sram_inv;
wire [0:3] sb_mux_size9_10_sram;
wire [0:3] sb_mux_size9_10_sram_inv;
wire [0:3] sb_mux_size9_11_sram;
wire [0:3] sb_mux_size9_11_sram_inv;
wire [0:3] sb_mux_size9_12_sram;
wire [0:3] sb_mux_size9_12_sram_inv;
wire [0:3] sb_mux_size9_13_sram;
wire [0:3] sb_mux_size9_13_sram_inv;
wire [0:3] sb_mux_size9_14_sram;
wire [0:3] sb_mux_size9_14_sram_inv;
wire [0:3] sb_mux_size9_15_sram;
wire [0:3] sb_mux_size9_15_sram_inv;
wire [0:3] sb_mux_size9_16_sram;
wire [0:3] sb_mux_size9_16_sram_inv;
wire [0:3] sb_mux_size9_17_sram;
wire [0:3] sb_mux_size9_17_sram_inv;
wire [0:3] sb_mux_size9_1_sram;
wire [0:3] sb_mux_size9_1_sram_inv;
wire [0:3] sb_mux_size9_2_sram;
wire [0:3] sb_mux_size9_2_sram_inv;
wire [0:3] sb_mux_size9_3_sram;
wire [0:3] sb_mux_size9_3_sram_inv;
wire [0:3] sb_mux_size9_4_sram;
wire [0:3] sb_mux_size9_4_sram_inv;
wire [0:3] sb_mux_size9_5_sram;
wire [0:3] sb_mux_size9_5_sram_inv;
wire [0:3] sb_mux_size9_6_sram;
wire [0:3] sb_mux_size9_6_sram_inv;
wire [0:3] sb_mux_size9_7_sram;
wire [0:3] sb_mux_size9_7_sram_inv;
wire [0:3] sb_mux_size9_8_sram;
wire [0:3] sb_mux_size9_8_sram_inv;
wire [0:3] sb_mux_size9_9_sram;
wire [0:3] sb_mux_size9_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[32] = chanx_right_in[32];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[33];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[34];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[35];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[36] = chanx_right_in[36];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[37];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[38];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[39];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[40] = chanx_right_in[40];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[41];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[42];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[43];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[44] = chanx_right_in[44];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[45];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[46];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[47];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[48];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[49];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[50];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[51];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[52] = chanx_right_in[52];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[53];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[54];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[55];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[56] = chanx_right_in[56];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[57];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[58];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[59];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[60] = chanx_right_in[60];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[61];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[62];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[63];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size11 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[1], chanx_right_in[6], chanx_right_in[26], bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[0], chanx_left_in[0], chanx_left_in[6], chanx_left_in[26]}),
		.sram(sb_mux_size11_0_sram[0:3]),
		.sram_inv(sb_mux_size11_0_sram_inv[0:3]),
		.out(chany_top_out[0]));

	sb_mux_size11 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[2], chanx_right_in[8], chanx_right_in[28], bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[1], chanx_left_in[8], chanx_left_in[28], chanx_left_in[31]}),
		.sram(sb_mux_size11_1_sram[0:3]),
		.sram_inv(sb_mux_size11_1_sram_inv[0:3]),
		.out(chany_top_out[1]));

	sb_mux_size11 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[9], chanx_right_in[16], bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[7], chanx_left_in[11], chanx_left_in[16]}),
		.sram(sb_mux_size11_2_sram[0:3]),
		.sram_inv(sb_mux_size11_2_sram_inv[0:3]),
		.out(chany_top_out[6]));

	sb_mux_size11 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[11], chanx_right_in[17], bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[9], chanx_left_in[9], chanx_left_in[17]}),
		.sram(sb_mux_size11_3_sram[0:3]),
		.sram_inv(sb_mux_size11_3_sram_inv[0:3]),
		.out(chany_top_out[8]));

	sb_mux_size11 mux_right_track_12 (
		.in({chany_top_in[5], chany_top_in[16], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_, chany_bottom_in[7], chany_bottom_in[16], chanx_left_in[7]}),
		.sram(sb_mux_size11_4_sram[0:3]),
		.sram_inv(sb_mux_size11_4_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	sb_mux_size11 mux_right_track_16 (
		.in({chany_top_in[7], chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_, chany_bottom_in[5], chany_bottom_in[17], chanx_left_in[9]}),
		.sram(sb_mux_size11_5_sram[0:3]),
		.sram_inv(sb_mux_size11_5_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	sb_mux_size11 mux_right_track_20 (
		.in({chany_top_in[9], chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_, chany_bottom_in[4], chany_bottom_in[18], chanx_left_in[11]}),
		.sram(sb_mux_size11_6_sram[0:3]),
		.sram_inv(sb_mux_size11_6_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	sb_mux_size11 mux_bottom_track_1 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_top_in[0], chanx_right_in[6], chanx_right_in[26:27], bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[1], chanx_left_in[6], chanx_left_in[26]}),
		.sram(sb_mux_size11_7_sram[0:3]),
		.sram_inv(sb_mux_size11_7_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	sb_mux_size11 mux_bottom_track_3 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_top_in[1], chanx_right_in[8], chanx_right_in[23], chanx_right_in[28], bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[2], chanx_left_in[8], chanx_left_in[28]}),
		.sram(sb_mux_size11_8_sram[0:3]),
		.sram_inv(sb_mux_size11_8_sram_inv[0:3]),
		.out(chany_bottom_out[1]));

	sb_mux_size11 mux_bottom_track_13 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_top_in[7], chanx_right_in[7], chanx_right_in[16], bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[9], chanx_left_in[16]}),
		.sram(sb_mux_size11_9_sram[0:3]),
		.sram_inv(sb_mux_size11_9_sram_inv[0:3]),
		.out(chany_bottom_out[6]));

	sb_mux_size11 mux_bottom_track_17 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_top_in[9], chanx_right_in[5], chanx_right_in[17], bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[11], chanx_left_in[17]}),
		.sram(sb_mux_size11_10_sram[0:3]),
		.sram_inv(sb_mux_size11_10_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	sb_mux_size11 mux_left_track_13 (
		.in({chany_top_in[11], chany_top_in[16], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_, chanx_right_in[7], chany_bottom_in[5], chany_bottom_in[16]}),
		.sram(sb_mux_size11_11_sram[0:3]),
		.sram_inv(sb_mux_size11_11_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	sb_mux_size11 mux_left_track_17 (
		.in({chany_top_in[9], chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_, chanx_right_in[9], chany_bottom_in[7], chany_bottom_in[17]}),
		.sram(sb_mux_size11_12_sram[0:3]),
		.sram_inv(sb_mux_size11_12_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	sb_mux_size11 mux_left_track_21 (
		.in({chany_top_in[7], chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_, chanx_right_in[11], chany_bottom_in[9], chany_bottom_in[18]}),
		.sram(sb_mux_size11_13_sram[0:3]),
		.sram_inv(sb_mux_size11_13_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_top_track_0 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[0:3]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[0:3]),
		.mem_out(sb_mux_size11_0_sram[0:3]),
		.mem_outb(sb_mux_size11_0_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_top_track_2 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[4:7]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[4:7]),
		.mem_out(sb_mux_size11_1_sram[0:3]),
		.mem_outb(sb_mux_size11_1_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_top_track_12 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[22:25]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[22:25]),
		.mem_out(sb_mux_size11_2_sram[0:3]),
		.mem_outb(sb_mux_size11_2_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_top_track_16 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[26:29]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[26:29]),
		.mem_out(sb_mux_size11_3_sram[0:3]),
		.mem_outb(sb_mux_size11_3_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_right_track_12 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[140:143]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[140:143]),
		.mem_out(sb_mux_size11_4_sram[0:3]),
		.mem_outb(sb_mux_size11_4_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_right_track_16 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[144:147]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[144:147]),
		.mem_out(sb_mux_size11_5_sram[0:3]),
		.mem_outb(sb_mux_size11_5_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_right_track_20 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[148:151]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[148:151]),
		.mem_out(sb_mux_size11_6_sram[0:3]),
		.mem_outb(sb_mux_size11_6_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_bottom_track_1 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[236:239]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[236:239]),
		.mem_out(sb_mux_size11_7_sram[0:3]),
		.mem_outb(sb_mux_size11_7_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_bottom_track_3 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[240:243]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[240:243]),
		.mem_out(sb_mux_size11_8_sram[0:3]),
		.mem_outb(sb_mux_size11_8_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_bottom_track_13 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[258:261]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[258:261]),
		.mem_out(sb_mux_size11_9_sram[0:3]),
		.mem_outb(sb_mux_size11_9_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_bottom_track_17 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[262:265]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[262:265]),
		.mem_out(sb_mux_size11_10_sram[0:3]),
		.mem_outb(sb_mux_size11_10_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_left_track_13 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[376:379]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[376:379]),
		.mem_out(sb_mux_size11_11_sram[0:3]),
		.mem_outb(sb_mux_size11_11_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_left_track_17 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[380:383]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[380:383]),
		.mem_out(sb_mux_size11_12_sram[0:3]),
		.mem_outb(sb_mux_size11_12_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_left_track_21 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[384:387]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[384:387]),
		.mem_out(sb_mux_size11_13_sram[0:3]),
		.mem_outb(sb_mux_size11_13_sram_inv[0:3]));

	sb_mux_size9 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_right_in[3], chanx_right_in[10], chanx_right_in[29], bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, chany_bottom_in[2], chanx_left_in[10], chanx_left_in[27], chanx_left_in[29]}),
		.sram(sb_mux_size9_0_sram[0:3]),
		.sram_inv(sb_mux_size9_0_sram_inv[0:3]),
		.out(chany_top_out[2]));

	sb_mux_size9 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[4], chanx_right_in[12], chanx_right_in[30], bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_bottom_in[3], chanx_left_in[12], chanx_left_in[23], chanx_left_in[30]}),
		.sram(sb_mux_size9_1_sram[0:3]),
		.sram_inv(sb_mux_size9_1_sram_inv[0:3]),
		.out(chany_top_out[3]));

	sb_mux_size9 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[15], chanx_right_in[18], bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[11], chanx_left_in[7], chanx_left_in[18]}),
		.sram(sb_mux_size9_2_sram[0:3]),
		.sram_inv(sb_mux_size9_2_sram_inv[0:3]),
		.out(chany_top_out[10]));

	sb_mux_size9 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[19:20], bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[15], chanx_left_in[5], chanx_left_in[20]}),
		.sram(sb_mux_size9_3_sram[0:3]),
		.sram_inv(sb_mux_size9_3_sram_inv[0:3]),
		.out(chany_top_out[12]));

	sb_mux_size9 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[21], chanx_right_in[23], bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[19], chanx_left_in[4], chanx_left_in[21]}),
		.sram(sb_mux_size9_4_sram[0:3]),
		.sram_inv(sb_mux_size9_4_sram_inv[0:3]),
		.out(chany_top_out[16]));

	sb_mux_size9 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[22], chanx_right_in[27], bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[23], chanx_left_in[3], chanx_left_in[22]}),
		.sram(sb_mux_size9_5_sram[0:3]),
		.sram_inv(sb_mux_size9_5_sram_inv[0:3]),
		.out(chany_top_out[20]));

	sb_mux_size9 mux_right_track_24 (
		.in({chany_top_in[11], chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_, chany_bottom_in[3], chany_bottom_in[20], chanx_left_in[15]}),
		.sram(sb_mux_size9_6_sram[0:3]),
		.sram_inv(sb_mux_size9_6_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	sb_mux_size9 mux_right_track_32 (
		.in({chany_top_in[15], chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_, chany_bottom_in[2], chany_bottom_in[21], chanx_left_in[19]}),
		.sram(sb_mux_size9_7_sram[0:3]),
		.sram_inv(sb_mux_size9_7_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	sb_mux_size9 mux_right_track_40 (
		.in({chany_top_in[19], chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_, chany_bottom_in[1], chany_bottom_in[22], chanx_left_in[23]}),
		.sram(sb_mux_size9_8_sram[0:3]),
		.sram_inv(sb_mux_size9_8_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	sb_mux_size9 mux_bottom_track_5 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, chany_top_in[2], chanx_right_in[10], chanx_right_in[19], chanx_right_in[29], bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_left_in[3], chanx_left_in[10], chanx_left_in[29]}),
		.sram(sb_mux_size9_9_sram[0:3]),
		.sram_inv(sb_mux_size9_9_sram_inv[0:3]),
		.out(chany_bottom_out[2]));

	sb_mux_size9 mux_bottom_track_7 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_top_in[3], chanx_right_in[12], chanx_right_in[15], chanx_right_in[30], bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_left_in[4], chanx_left_in[12], chanx_left_in[30]}),
		.sram(sb_mux_size9_10_sram[0:3]),
		.sram_inv(sb_mux_size9_10_sram_inv[0:3]),
		.out(chany_bottom_out[3]));

	sb_mux_size9 mux_bottom_track_21 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_top_in[11], chanx_right_in[4], chanx_right_in[18], bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[15], chanx_left_in[18]}),
		.sram(sb_mux_size9_11_sram[0:3]),
		.sram_inv(sb_mux_size9_11_sram_inv[0:3]),
		.out(chany_bottom_out[10]));

	sb_mux_size9 mux_bottom_track_25 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_top_in[15], chanx_right_in[3], chanx_right_in[20], bottom_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[19:20]}),
		.sram(sb_mux_size9_12_sram[0:3]),
		.sram_inv(sb_mux_size9_12_sram_inv[0:3]),
		.out(chany_bottom_out[12]));

	sb_mux_size9 mux_bottom_track_33 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_top_in[19], chanx_right_in[2], chanx_right_in[21], bottom_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[21], chanx_left_in[23]}),
		.sram(sb_mux_size9_13_sram[0:3]),
		.sram_inv(sb_mux_size9_13_sram_inv[0:3]),
		.out(chany_bottom_out[16]));

	sb_mux_size9 mux_bottom_track_41 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_top_in[23], chanx_right_in[1], chanx_right_in[22], bottom_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[22], chanx_left_in[27]}),
		.sram(sb_mux_size9_14_sram[0:3]),
		.sram_inv(sb_mux_size9_14_sram_inv[0:3]),
		.out(chany_bottom_out[20]));

	sb_mux_size9 mux_left_track_25 (
		.in({chany_top_in[5], chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_, chanx_right_in[15], chany_bottom_in[11], chany_bottom_in[20]}),
		.sram(sb_mux_size9_15_sram[0:3]),
		.sram_inv(sb_mux_size9_15_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	sb_mux_size9 mux_left_track_33 (
		.in({chany_top_in[4], chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_, chanx_right_in[19], chany_bottom_in[15], chany_bottom_in[21]}),
		.sram(sb_mux_size9_16_sram[0:3]),
		.sram_inv(sb_mux_size9_16_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	sb_mux_size9 mux_left_track_41 (
		.in({chany_top_in[3], chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_, chanx_right_in[23], chany_bottom_in[19], chany_bottom_in[22]}),
		.sram(sb_mux_size9_17_sram[0:3]),
		.sram_inv(sb_mux_size9_17_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_4 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[8:11]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[8:11]),
		.mem_out(sb_mux_size9_0_sram[0:3]),
		.mem_outb(sb_mux_size9_0_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_6 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[12:15]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[12:15]),
		.mem_out(sb_mux_size9_1_sram[0:3]),
		.mem_outb(sb_mux_size9_1_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_20 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[30:33]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[30:33]),
		.mem_out(sb_mux_size9_2_sram[0:3]),
		.mem_outb(sb_mux_size9_2_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_24 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[34:37]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[34:37]),
		.mem_out(sb_mux_size9_3_sram[0:3]),
		.mem_outb(sb_mux_size9_3_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_32 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[38:41]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[38:41]),
		.mem_out(sb_mux_size9_4_sram[0:3]),
		.mem_outb(sb_mux_size9_4_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_40 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[42:45]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[42:45]),
		.mem_out(sb_mux_size9_5_sram[0:3]),
		.mem_outb(sb_mux_size9_5_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_24 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[152:155]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[152:155]),
		.mem_out(sb_mux_size9_6_sram[0:3]),
		.mem_outb(sb_mux_size9_6_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_32 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[156:159]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[156:159]),
		.mem_out(sb_mux_size9_7_sram[0:3]),
		.mem_outb(sb_mux_size9_7_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_40 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[160:163]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[160:163]),
		.mem_out(sb_mux_size9_8_sram[0:3]),
		.mem_outb(sb_mux_size9_8_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_bottom_track_5 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[244:247]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[244:247]),
		.mem_out(sb_mux_size9_9_sram[0:3]),
		.mem_outb(sb_mux_size9_9_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_bottom_track_7 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[248:251]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[248:251]),
		.mem_out(sb_mux_size9_10_sram[0:3]),
		.mem_outb(sb_mux_size9_10_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_bottom_track_21 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[266:269]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[266:269]),
		.mem_out(sb_mux_size9_11_sram[0:3]),
		.mem_outb(sb_mux_size9_11_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_bottom_track_25 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[270:273]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[270:273]),
		.mem_out(sb_mux_size9_12_sram[0:3]),
		.mem_outb(sb_mux_size9_12_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_bottom_track_33 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[274:277]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[274:277]),
		.mem_out(sb_mux_size9_13_sram[0:3]),
		.mem_outb(sb_mux_size9_13_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_bottom_track_41 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[278:281]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[278:281]),
		.mem_out(sb_mux_size9_14_sram[0:3]),
		.mem_outb(sb_mux_size9_14_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_25 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[388:391]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[388:391]),
		.mem_out(sb_mux_size9_15_sram[0:3]),
		.mem_outb(sb_mux_size9_15_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_33 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[392:395]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[392:395]),
		.mem_out(sb_mux_size9_16_sram[0:3]),
		.mem_outb(sb_mux_size9_16_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_41 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[396:399]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[396:399]),
		.mem_out(sb_mux_size9_17_sram[0:3]),
		.mem_outb(sb_mux_size9_17_sram_inv[0:3]));

	sb_mux_size7 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[5], chanx_right_in[13], bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_bottom_in[4], chanx_left_in[13], chanx_left_in[19]}),
		.sram(sb_mux_size7_0_sram[0:2]),
		.sram_inv(sb_mux_size7_0_sram_inv[0:2]),
		.out(chany_top_out[4]));

	sb_mux_size7 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[7], chanx_right_in[14], bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[5], chanx_left_in[14:15]}),
		.sram(sb_mux_size7_1_sram[0:2]),
		.sram_inv(sb_mux_size7_1_sram_inv[0:2]),
		.out(chany_top_out[5]));

	sb_mux_size7 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[24], chanx_right_in[31], bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_bottom_in[27], chanx_left_in[2], chanx_left_in[24]}),
		.sram(sb_mux_size7_2_sram[0:2]),
		.sram_inv(sb_mux_size7_2_sram_inv[0:2]),
		.out(chany_top_out[24]));

	sb_mux_size7 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[0], chanx_right_in[25], bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_bottom_in[31], chanx_left_in[1], chanx_left_in[25]}),
		.sram(sb_mux_size7_3_sram[0:2]),
		.sram_inv(sb_mux_size7_3_sram_inv[0:2]),
		.out(chany_top_out[28]));

	sb_mux_size7 mux_bottom_track_9 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_top_in[4], chanx_right_in[11], chanx_right_in[13], bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_left_in[5], chanx_left_in[13]}),
		.sram(sb_mux_size7_4_sram[0:2]),
		.sram_inv(sb_mux_size7_4_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	sb_mux_size7 mux_bottom_track_11 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_top_in[5], chanx_right_in[9], chanx_right_in[14], bottom_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[7], chanx_left_in[14]}),
		.sram(sb_mux_size7_5_sram[0:2]),
		.sram_inv(sb_mux_size7_5_sram_inv[0:2]),
		.out(chany_bottom_out[5]));

	sb_mux_size7 mux_bottom_track_49 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_top_in[27], chanx_right_in[0], chanx_right_in[24], bottom_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_left_in[24], chanx_left_in[31]}),
		.sram(sb_mux_size7_6_sram[0:2]),
		.sram_inv(sb_mux_size7_6_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	sb_mux_size7 mux_bottom_track_57 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_top_in[31], chanx_right_in[25], chanx_right_in[31], bottom_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_left_in[0], chanx_left_in[25]}),
		.sram(sb_mux_size7_7_sram[0:2]),
		.sram_inv(sb_mux_size7_7_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_8 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[16:18]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[16:18]),
		.mem_out(sb_mux_size7_0_sram[0:2]),
		.mem_outb(sb_mux_size7_0_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_10 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[19:21]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[19:21]),
		.mem_out(sb_mux_size7_1_sram[0:2]),
		.mem_outb(sb_mux_size7_1_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_48 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[46:48]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[46:48]),
		.mem_out(sb_mux_size7_2_sram[0:2]),
		.mem_outb(sb_mux_size7_2_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_56 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[49:51]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[49:51]),
		.mem_out(sb_mux_size7_3_sram[0:2]),
		.mem_outb(sb_mux_size7_3_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_9 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[252:254]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[252:254]),
		.mem_out(sb_mux_size7_4_sram[0:2]),
		.mem_outb(sb_mux_size7_4_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_11 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[255:257]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[255:257]),
		.mem_out(sb_mux_size7_5_sram[0:2]),
		.mem_outb(sb_mux_size7_5_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_49 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[282:284]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[282:284]),
		.mem_out(sb_mux_size7_6_sram[0:2]),
		.mem_outb(sb_mux_size7_6_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_57 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[285:287]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[285:287]),
		.mem_out(sb_mux_size7_7_sram[0:2]),
		.mem_outb(sb_mux_size7_7_sram_inv[0:2]));

	clk_mux_size3 mux_top_track_64 (
		.in({chanx_right_in[32], chany_bottom_in[32], chanx_left_in[32]}),
		.sram(clk_mux_size3_0_sram[0:1]),
		.sram_inv(clk_mux_size3_0_sram_inv[0:1]),
		.out(chany_top_out[32]));

	clk_mux_size3 mux_top_track_66 (
		.in({chanx_right_in[33], chany_bottom_in[33], chanx_left_in[33]}),
		.sram(clk_mux_size3_1_sram[0:1]),
		.sram_inv(clk_mux_size3_1_sram_inv[0:1]),
		.out(chany_top_out[33]));

	clk_mux_size3 mux_top_track_68 (
		.in({chanx_right_in[34], chany_bottom_in[34], chanx_left_in[34]}),
		.sram(clk_mux_size3_2_sram[0:1]),
		.sram_inv(clk_mux_size3_2_sram_inv[0:1]),
		.out(chany_top_out[34]));

	clk_mux_size3 mux_top_track_70 (
		.in({chanx_right_in[35], chany_bottom_in[35], chanx_left_in[35]}),
		.sram(clk_mux_size3_3_sram[0:1]),
		.sram_inv(clk_mux_size3_3_sram_inv[0:1]),
		.out(chany_top_out[35]));

	clk_mux_size3 mux_top_track_72 (
		.in({chanx_right_in[36], chany_bottom_in[36], chanx_left_in[36]}),
		.sram(clk_mux_size3_4_sram[0:1]),
		.sram_inv(clk_mux_size3_4_sram_inv[0:1]),
		.out(chany_top_out[36]));

	clk_mux_size3 mux_top_track_74 (
		.in({chanx_right_in[37], chany_bottom_in[37], chanx_left_in[37]}),
		.sram(clk_mux_size3_5_sram[0:1]),
		.sram_inv(clk_mux_size3_5_sram_inv[0:1]),
		.out(chany_top_out[37]));

	clk_mux_size3 mux_top_track_76 (
		.in({chanx_right_in[38], chany_bottom_in[38], chanx_left_in[38]}),
		.sram(clk_mux_size3_6_sram[0:1]),
		.sram_inv(clk_mux_size3_6_sram_inv[0:1]),
		.out(chany_top_out[38]));

	clk_mux_size3 mux_top_track_78 (
		.in({chanx_right_in[39], chany_bottom_in[39], chanx_left_in[39]}),
		.sram(clk_mux_size3_7_sram[0:1]),
		.sram_inv(clk_mux_size3_7_sram_inv[0:1]),
		.out(chany_top_out[39]));

	clk_mux_size3 mux_top_track_80 (
		.in({chanx_right_in[40], chany_bottom_in[40], chanx_left_in[40]}),
		.sram(clk_mux_size3_8_sram[0:1]),
		.sram_inv(clk_mux_size3_8_sram_inv[0:1]),
		.out(chany_top_out[40]));

	clk_mux_size3 mux_top_track_82 (
		.in({chanx_right_in[41], chany_bottom_in[41], chanx_left_in[41]}),
		.sram(clk_mux_size3_9_sram[0:1]),
		.sram_inv(clk_mux_size3_9_sram_inv[0:1]),
		.out(chany_top_out[41]));

	clk_mux_size3 mux_top_track_84 (
		.in({chanx_right_in[42], chany_bottom_in[42], chanx_left_in[42]}),
		.sram(clk_mux_size3_10_sram[0:1]),
		.sram_inv(clk_mux_size3_10_sram_inv[0:1]),
		.out(chany_top_out[42]));

	clk_mux_size3 mux_top_track_86 (
		.in({chanx_right_in[43], chany_bottom_in[43], chanx_left_in[43]}),
		.sram(clk_mux_size3_11_sram[0:1]),
		.sram_inv(clk_mux_size3_11_sram_inv[0:1]),
		.out(chany_top_out[43]));

	clk_mux_size3 mux_top_track_88 (
		.in({chanx_right_in[44], chany_bottom_in[44], chanx_left_in[44]}),
		.sram(clk_mux_size3_12_sram[0:1]),
		.sram_inv(clk_mux_size3_12_sram_inv[0:1]),
		.out(chany_top_out[44]));

	clk_mux_size3 mux_top_track_90 (
		.in({chanx_right_in[45], chany_bottom_in[45], chanx_left_in[45]}),
		.sram(clk_mux_size3_13_sram[0:1]),
		.sram_inv(clk_mux_size3_13_sram_inv[0:1]),
		.out(chany_top_out[45]));

	clk_mux_size3 mux_top_track_92 (
		.in({chanx_right_in[46], chany_bottom_in[46], chanx_left_in[46]}),
		.sram(clk_mux_size3_14_sram[0:1]),
		.sram_inv(clk_mux_size3_14_sram_inv[0:1]),
		.out(chany_top_out[46]));

	clk_mux_size3 mux_top_track_94 (
		.in({chanx_right_in[47], chany_bottom_in[47], chanx_left_in[47]}),
		.sram(clk_mux_size3_15_sram[0:1]),
		.sram_inv(clk_mux_size3_15_sram_inv[0:1]),
		.out(chany_top_out[47]));

	clk_mux_size3 mux_top_track_96 (
		.in({chanx_right_in[48], chany_bottom_in[48], chanx_left_in[48]}),
		.sram(clk_mux_size3_16_sram[0:1]),
		.sram_inv(clk_mux_size3_16_sram_inv[0:1]),
		.out(chany_top_out[48]));

	clk_mux_size3 mux_top_track_98 (
		.in({chanx_right_in[49], chany_bottom_in[49], chanx_left_in[49]}),
		.sram(clk_mux_size3_17_sram[0:1]),
		.sram_inv(clk_mux_size3_17_sram_inv[0:1]),
		.out(chany_top_out[49]));

	clk_mux_size3 mux_top_track_100 (
		.in({chanx_right_in[50], chany_bottom_in[50], chanx_left_in[50]}),
		.sram(clk_mux_size3_18_sram[0:1]),
		.sram_inv(clk_mux_size3_18_sram_inv[0:1]),
		.out(chany_top_out[50]));

	clk_mux_size3 mux_top_track_102 (
		.in({chanx_right_in[51], chany_bottom_in[51], chanx_left_in[51]}),
		.sram(clk_mux_size3_19_sram[0:1]),
		.sram_inv(clk_mux_size3_19_sram_inv[0:1]),
		.out(chany_top_out[51]));

	clk_mux_size3 mux_top_track_104 (
		.in({chanx_right_in[52], chany_bottom_in[52], chanx_left_in[52]}),
		.sram(clk_mux_size3_20_sram[0:1]),
		.sram_inv(clk_mux_size3_20_sram_inv[0:1]),
		.out(chany_top_out[52]));

	clk_mux_size3 mux_top_track_106 (
		.in({chanx_right_in[53], chany_bottom_in[53], chanx_left_in[53]}),
		.sram(clk_mux_size3_21_sram[0:1]),
		.sram_inv(clk_mux_size3_21_sram_inv[0:1]),
		.out(chany_top_out[53]));

	clk_mux_size3 mux_top_track_108 (
		.in({chanx_right_in[54], chany_bottom_in[54], chanx_left_in[54]}),
		.sram(clk_mux_size3_22_sram[0:1]),
		.sram_inv(clk_mux_size3_22_sram_inv[0:1]),
		.out(chany_top_out[54]));

	clk_mux_size3 mux_top_track_110 (
		.in({chanx_right_in[55], chany_bottom_in[55], chanx_left_in[55]}),
		.sram(clk_mux_size3_23_sram[0:1]),
		.sram_inv(clk_mux_size3_23_sram_inv[0:1]),
		.out(chany_top_out[55]));

	clk_mux_size3 mux_top_track_112 (
		.in({chanx_right_in[56], chany_bottom_in[56], chanx_left_in[56]}),
		.sram(clk_mux_size3_24_sram[0:1]),
		.sram_inv(clk_mux_size3_24_sram_inv[0:1]),
		.out(chany_top_out[56]));

	clk_mux_size3 mux_top_track_114 (
		.in({chanx_right_in[57], chany_bottom_in[57], chanx_left_in[57]}),
		.sram(clk_mux_size3_25_sram[0:1]),
		.sram_inv(clk_mux_size3_25_sram_inv[0:1]),
		.out(chany_top_out[57]));

	clk_mux_size3 mux_top_track_116 (
		.in({chanx_right_in[58], chany_bottom_in[58], chanx_left_in[58]}),
		.sram(clk_mux_size3_26_sram[0:1]),
		.sram_inv(clk_mux_size3_26_sram_inv[0:1]),
		.out(chany_top_out[58]));

	clk_mux_size3 mux_top_track_118 (
		.in({chanx_right_in[59], chany_bottom_in[59], chanx_left_in[59]}),
		.sram(clk_mux_size3_27_sram[0:1]),
		.sram_inv(clk_mux_size3_27_sram_inv[0:1]),
		.out(chany_top_out[59]));

	clk_mux_size3 mux_top_track_120 (
		.in({chanx_right_in[60], chany_bottom_in[60], chanx_left_in[60]}),
		.sram(clk_mux_size3_28_sram[0:1]),
		.sram_inv(clk_mux_size3_28_sram_inv[0:1]),
		.out(chany_top_out[60]));

	clk_mux_size3 mux_top_track_122 (
		.in({chanx_right_in[61], chany_bottom_in[61], chanx_left_in[61]}),
		.sram(clk_mux_size3_29_sram[0:1]),
		.sram_inv(clk_mux_size3_29_sram_inv[0:1]),
		.out(chany_top_out[61]));

	clk_mux_size3 mux_top_track_124 (
		.in({chanx_right_in[62], chany_bottom_in[62], chanx_left_in[62]}),
		.sram(clk_mux_size3_30_sram[0:1]),
		.sram_inv(clk_mux_size3_30_sram_inv[0:1]),
		.out(chany_top_out[62]));

	clk_mux_size3 mux_top_track_126 (
		.in({chanx_right_in[63], chany_bottom_in[63], chanx_left_in[63]}),
		.sram(clk_mux_size3_31_sram[0:1]),
		.sram_inv(clk_mux_size3_31_sram_inv[0:1]),
		.out(chany_top_out[63]));

	clk_mux_size3 mux_right_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_out_0_, chanx_left_in[32]}),
		.sram(clk_mux_size3_32_sram[0:1]),
		.sram_inv(clk_mux_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	clk_mux_size3 mux_right_track_66 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_out_0_, chanx_left_in[33]}),
		.sram(clk_mux_size3_33_sram[0:1]),
		.sram_inv(clk_mux_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	clk_mux_size3 mux_right_track_68 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_out_0_, chanx_left_in[34]}),
		.sram(clk_mux_size3_34_sram[0:1]),
		.sram_inv(clk_mux_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	clk_mux_size3 mux_right_track_70 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_out_0_, chanx_left_in[35]}),
		.sram(clk_mux_size3_35_sram[0:1]),
		.sram_inv(clk_mux_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	clk_mux_size3 mux_right_track_72 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_out_0_, chanx_left_in[36]}),
		.sram(clk_mux_size3_36_sram[0:1]),
		.sram_inv(clk_mux_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	clk_mux_size3 mux_right_track_74 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_out_0_, chanx_left_in[37]}),
		.sram(clk_mux_size3_37_sram[0:1]),
		.sram_inv(clk_mux_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	clk_mux_size3 mux_right_track_76 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_out_0_, chanx_left_in[38]}),
		.sram(clk_mux_size3_38_sram[0:1]),
		.sram_inv(clk_mux_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	clk_mux_size3 mux_right_track_78 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_out_0_, chanx_left_in[39]}),
		.sram(clk_mux_size3_39_sram[0:1]),
		.sram_inv(clk_mux_size3_39_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	clk_mux_size3 mux_right_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_8__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_8__pin_out_0_, chanx_left_in[40]}),
		.sram(clk_mux_size3_40_sram[0:1]),
		.sram_inv(clk_mux_size3_40_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	clk_mux_size3 mux_right_track_82 (
		.in({top_right_grid_left_width_0_height_0_subtile_9__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_9__pin_out_0_, chanx_left_in[41]}),
		.sram(clk_mux_size3_41_sram[0:1]),
		.sram_inv(clk_mux_size3_41_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	clk_mux_size3 mux_right_track_84 (
		.in({top_right_grid_left_width_0_height_0_subtile_10__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_10__pin_out_0_, chanx_left_in[42]}),
		.sram(clk_mux_size3_42_sram[0:1]),
		.sram_inv(clk_mux_size3_42_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	clk_mux_size3 mux_right_track_86 (
		.in({top_right_grid_left_width_0_height_0_subtile_11__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_11__pin_out_0_, chanx_left_in[43]}),
		.sram(clk_mux_size3_43_sram[0:1]),
		.sram_inv(clk_mux_size3_43_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	clk_mux_size3 mux_right_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_12__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_12__pin_out_0_, chanx_left_in[44]}),
		.sram(clk_mux_size3_44_sram[0:1]),
		.sram_inv(clk_mux_size3_44_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	clk_mux_size3 mux_right_track_90 (
		.in({top_right_grid_left_width_0_height_0_subtile_13__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_13__pin_out_0_, chanx_left_in[45]}),
		.sram(clk_mux_size3_45_sram[0:1]),
		.sram_inv(clk_mux_size3_45_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	clk_mux_size3 mux_right_track_92 (
		.in({top_right_grid_left_width_0_height_0_subtile_14__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_14__pin_out_0_, chanx_left_in[46]}),
		.sram(clk_mux_size3_46_sram[0:1]),
		.sram_inv(clk_mux_size3_46_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	clk_mux_size3 mux_right_track_94 (
		.in({top_right_grid_left_width_0_height_0_subtile_15__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_15__pin_out_0_, chanx_left_in[47]}),
		.sram(clk_mux_size3_47_sram[0:1]),
		.sram_inv(clk_mux_size3_47_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	clk_mux_size3 mux_right_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_16__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_16__pin_out_0_, chanx_left_in[48]}),
		.sram(clk_mux_size3_48_sram[0:1]),
		.sram_inv(clk_mux_size3_48_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	clk_mux_size3 mux_right_track_98 (
		.in({top_right_grid_left_width_0_height_0_subtile_17__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_17__pin_out_0_, chanx_left_in[49]}),
		.sram(clk_mux_size3_49_sram[0:1]),
		.sram_inv(clk_mux_size3_49_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	clk_mux_size3 mux_right_track_100 (
		.in({top_right_grid_left_width_0_height_0_subtile_18__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_18__pin_out_0_, chanx_left_in[50]}),
		.sram(clk_mux_size3_50_sram[0:1]),
		.sram_inv(clk_mux_size3_50_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	clk_mux_size3 mux_right_track_102 (
		.in({top_right_grid_left_width_0_height_0_subtile_19__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_19__pin_out_0_, chanx_left_in[51]}),
		.sram(clk_mux_size3_51_sram[0:1]),
		.sram_inv(clk_mux_size3_51_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	clk_mux_size3 mux_right_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_8__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_8__pin_out_0_, chanx_left_in[52]}),
		.sram(clk_mux_size3_52_sram[0:1]),
		.sram_inv(clk_mux_size3_52_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	clk_mux_size3 mux_right_track_106 (
		.in({top_right_grid_left_width_0_height_0_subtile_9__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_9__pin_out_0_, chanx_left_in[53]}),
		.sram(clk_mux_size3_53_sram[0:1]),
		.sram_inv(clk_mux_size3_53_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	clk_mux_size3 mux_right_track_108 (
		.in({top_right_grid_left_width_0_height_0_subtile_10__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_10__pin_out_0_, chanx_left_in[54]}),
		.sram(clk_mux_size3_54_sram[0:1]),
		.sram_inv(clk_mux_size3_54_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	clk_mux_size3 mux_right_track_110 (
		.in({top_right_grid_left_width_0_height_0_subtile_11__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_11__pin_out_0_, chanx_left_in[55]}),
		.sram(clk_mux_size3_55_sram[0:1]),
		.sram_inv(clk_mux_size3_55_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	clk_mux_size3 mux_right_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_12__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_12__pin_out_0_, chanx_left_in[56]}),
		.sram(clk_mux_size3_56_sram[0:1]),
		.sram_inv(clk_mux_size3_56_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	clk_mux_size3 mux_right_track_114 (
		.in({top_right_grid_left_width_0_height_0_subtile_13__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_13__pin_out_0_, chanx_left_in[57]}),
		.sram(clk_mux_size3_57_sram[0:1]),
		.sram_inv(clk_mux_size3_57_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	clk_mux_size3 mux_right_track_116 (
		.in({top_right_grid_left_width_0_height_0_subtile_14__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_14__pin_out_0_, chanx_left_in[58]}),
		.sram(clk_mux_size3_58_sram[0:1]),
		.sram_inv(clk_mux_size3_58_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	clk_mux_size3 mux_right_track_118 (
		.in({top_right_grid_left_width_0_height_0_subtile_15__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_15__pin_out_0_, chanx_left_in[59]}),
		.sram(clk_mux_size3_59_sram[0:1]),
		.sram_inv(clk_mux_size3_59_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	clk_mux_size3 mux_right_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_16__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_16__pin_out_0_, chanx_left_in[60]}),
		.sram(clk_mux_size3_60_sram[0:1]),
		.sram_inv(clk_mux_size3_60_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	clk_mux_size3 mux_right_track_122 (
		.in({top_right_grid_left_width_0_height_0_subtile_17__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_17__pin_out_0_, chanx_left_in[61]}),
		.sram(clk_mux_size3_61_sram[0:1]),
		.sram_inv(clk_mux_size3_61_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	clk_mux_size3 mux_right_track_124 (
		.in({top_right_grid_left_width_0_height_0_subtile_18__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_18__pin_out_0_, chanx_left_in[62]}),
		.sram(clk_mux_size3_62_sram[0:1]),
		.sram_inv(clk_mux_size3_62_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	clk_mux_size3 mux_right_track_126 (
		.in({top_right_grid_left_width_0_height_0_subtile_19__pin_out_0_, bottom_right_grid_left_width_0_height_0_subtile_19__pin_out_0_, chanx_left_in[63]}),
		.sram(clk_mux_size3_63_sram[0:1]),
		.sram_inv(clk_mux_size3_63_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	clk_mux_size3 mux_bottom_track_65 (
		.in({chany_top_in[32], chanx_right_in[32], chanx_left_in[32]}),
		.sram(clk_mux_size3_64_sram[0:1]),
		.sram_inv(clk_mux_size3_64_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	clk_mux_size3 mux_bottom_track_67 (
		.in({chany_top_in[33], chanx_right_in[33], chanx_left_in[33]}),
		.sram(clk_mux_size3_65_sram[0:1]),
		.sram_inv(clk_mux_size3_65_sram_inv[0:1]),
		.out(chany_bottom_out[33]));

	clk_mux_size3 mux_bottom_track_69 (
		.in({chany_top_in[34], chanx_right_in[34], chanx_left_in[34]}),
		.sram(clk_mux_size3_66_sram[0:1]),
		.sram_inv(clk_mux_size3_66_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	clk_mux_size3 mux_bottom_track_71 (
		.in({chany_top_in[35], chanx_right_in[35], chanx_left_in[35]}),
		.sram(clk_mux_size3_67_sram[0:1]),
		.sram_inv(clk_mux_size3_67_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	clk_mux_size3 mux_bottom_track_73 (
		.in({chany_top_in[36], chanx_right_in[36], chanx_left_in[36]}),
		.sram(clk_mux_size3_68_sram[0:1]),
		.sram_inv(clk_mux_size3_68_sram_inv[0:1]),
		.out(chany_bottom_out[36]));

	clk_mux_size3 mux_bottom_track_75 (
		.in({chany_top_in[37], chanx_right_in[37], chanx_left_in[37]}),
		.sram(clk_mux_size3_69_sram[0:1]),
		.sram_inv(clk_mux_size3_69_sram_inv[0:1]),
		.out(chany_bottom_out[37]));

	clk_mux_size3 mux_bottom_track_77 (
		.in({chany_top_in[38], chanx_right_in[38], chanx_left_in[38]}),
		.sram(clk_mux_size3_70_sram[0:1]),
		.sram_inv(clk_mux_size3_70_sram_inv[0:1]),
		.out(chany_bottom_out[38]));

	clk_mux_size3 mux_bottom_track_79 (
		.in({chany_top_in[39], chanx_right_in[39], chanx_left_in[39]}),
		.sram(clk_mux_size3_71_sram[0:1]),
		.sram_inv(clk_mux_size3_71_sram_inv[0:1]),
		.out(chany_bottom_out[39]));

	clk_mux_size3 mux_bottom_track_81 (
		.in({chany_top_in[40], chanx_right_in[40], chanx_left_in[40]}),
		.sram(clk_mux_size3_72_sram[0:1]),
		.sram_inv(clk_mux_size3_72_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	clk_mux_size3 mux_bottom_track_83 (
		.in({chany_top_in[41], chanx_right_in[41], chanx_left_in[41]}),
		.sram(clk_mux_size3_73_sram[0:1]),
		.sram_inv(clk_mux_size3_73_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	clk_mux_size3 mux_bottom_track_85 (
		.in({chany_top_in[42], chanx_right_in[42], chanx_left_in[42]}),
		.sram(clk_mux_size3_74_sram[0:1]),
		.sram_inv(clk_mux_size3_74_sram_inv[0:1]),
		.out(chany_bottom_out[42]));

	clk_mux_size3 mux_bottom_track_87 (
		.in({chany_top_in[43], chanx_right_in[43], chanx_left_in[43]}),
		.sram(clk_mux_size3_75_sram[0:1]),
		.sram_inv(clk_mux_size3_75_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	clk_mux_size3 mux_bottom_track_89 (
		.in({chany_top_in[44], chanx_right_in[44], chanx_left_in[44]}),
		.sram(clk_mux_size3_76_sram[0:1]),
		.sram_inv(clk_mux_size3_76_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	clk_mux_size3 mux_bottom_track_91 (
		.in({chany_top_in[45], chanx_right_in[45], chanx_left_in[45]}),
		.sram(clk_mux_size3_77_sram[0:1]),
		.sram_inv(clk_mux_size3_77_sram_inv[0:1]),
		.out(chany_bottom_out[45]));

	clk_mux_size3 mux_bottom_track_93 (
		.in({chany_top_in[46], chanx_right_in[46], chanx_left_in[46]}),
		.sram(clk_mux_size3_78_sram[0:1]),
		.sram_inv(clk_mux_size3_78_sram_inv[0:1]),
		.out(chany_bottom_out[46]));

	clk_mux_size3 mux_bottom_track_95 (
		.in({chany_top_in[47], chanx_right_in[47], chanx_left_in[47]}),
		.sram(clk_mux_size3_79_sram[0:1]),
		.sram_inv(clk_mux_size3_79_sram_inv[0:1]),
		.out(chany_bottom_out[47]));

	clk_mux_size3 mux_bottom_track_97 (
		.in({chany_top_in[48], chanx_right_in[48], chanx_left_in[48]}),
		.sram(clk_mux_size3_80_sram[0:1]),
		.sram_inv(clk_mux_size3_80_sram_inv[0:1]),
		.out(chany_bottom_out[48]));

	clk_mux_size3 mux_bottom_track_99 (
		.in({chany_top_in[49], chanx_right_in[49], chanx_left_in[49]}),
		.sram(clk_mux_size3_81_sram[0:1]),
		.sram_inv(clk_mux_size3_81_sram_inv[0:1]),
		.out(chany_bottom_out[49]));

	clk_mux_size3 mux_bottom_track_101 (
		.in({chany_top_in[50], chanx_right_in[50], chanx_left_in[50]}),
		.sram(clk_mux_size3_82_sram[0:1]),
		.sram_inv(clk_mux_size3_82_sram_inv[0:1]),
		.out(chany_bottom_out[50]));

	clk_mux_size3 mux_bottom_track_103 (
		.in({chany_top_in[51], chanx_right_in[51], chanx_left_in[51]}),
		.sram(clk_mux_size3_83_sram[0:1]),
		.sram_inv(clk_mux_size3_83_sram_inv[0:1]),
		.out(chany_bottom_out[51]));

	clk_mux_size3 mux_bottom_track_105 (
		.in({chany_top_in[52], chanx_right_in[52], chanx_left_in[52]}),
		.sram(clk_mux_size3_84_sram[0:1]),
		.sram_inv(clk_mux_size3_84_sram_inv[0:1]),
		.out(chany_bottom_out[52]));

	clk_mux_size3 mux_bottom_track_107 (
		.in({chany_top_in[53], chanx_right_in[53], chanx_left_in[53]}),
		.sram(clk_mux_size3_85_sram[0:1]),
		.sram_inv(clk_mux_size3_85_sram_inv[0:1]),
		.out(chany_bottom_out[53]));

	clk_mux_size3 mux_bottom_track_109 (
		.in({chany_top_in[54], chanx_right_in[54], chanx_left_in[54]}),
		.sram(clk_mux_size3_86_sram[0:1]),
		.sram_inv(clk_mux_size3_86_sram_inv[0:1]),
		.out(chany_bottom_out[54]));

	clk_mux_size3 mux_bottom_track_111 (
		.in({chany_top_in[55], chanx_right_in[55], chanx_left_in[55]}),
		.sram(clk_mux_size3_87_sram[0:1]),
		.sram_inv(clk_mux_size3_87_sram_inv[0:1]),
		.out(chany_bottom_out[55]));

	clk_mux_size3 mux_bottom_track_113 (
		.in({chany_top_in[56], chanx_right_in[56], chanx_left_in[56]}),
		.sram(clk_mux_size3_88_sram[0:1]),
		.sram_inv(clk_mux_size3_88_sram_inv[0:1]),
		.out(chany_bottom_out[56]));

	clk_mux_size3 mux_bottom_track_115 (
		.in({chany_top_in[57], chanx_right_in[57], chanx_left_in[57]}),
		.sram(clk_mux_size3_89_sram[0:1]),
		.sram_inv(clk_mux_size3_89_sram_inv[0:1]),
		.out(chany_bottom_out[57]));

	clk_mux_size3 mux_bottom_track_117 (
		.in({chany_top_in[58], chanx_right_in[58], chanx_left_in[58]}),
		.sram(clk_mux_size3_90_sram[0:1]),
		.sram_inv(clk_mux_size3_90_sram_inv[0:1]),
		.out(chany_bottom_out[58]));

	clk_mux_size3 mux_bottom_track_119 (
		.in({chany_top_in[59], chanx_right_in[59], chanx_left_in[59]}),
		.sram(clk_mux_size3_91_sram[0:1]),
		.sram_inv(clk_mux_size3_91_sram_inv[0:1]),
		.out(chany_bottom_out[59]));

	clk_mux_size3 mux_bottom_track_121 (
		.in({chany_top_in[60], chanx_right_in[60], chanx_left_in[60]}),
		.sram(clk_mux_size3_92_sram[0:1]),
		.sram_inv(clk_mux_size3_92_sram_inv[0:1]),
		.out(chany_bottom_out[60]));

	clk_mux_size3 mux_bottom_track_123 (
		.in({chany_top_in[61], chanx_right_in[61], chanx_left_in[61]}),
		.sram(clk_mux_size3_93_sram[0:1]),
		.sram_inv(clk_mux_size3_93_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	clk_mux_size3 mux_bottom_track_125 (
		.in({chany_top_in[62], chanx_right_in[62], chanx_left_in[62]}),
		.sram(clk_mux_size3_94_sram[0:1]),
		.sram_inv(clk_mux_size3_94_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	clk_mux_size3 mux_bottom_track_127 (
		.in({chany_top_in[63], chanx_right_in[63], chanx_left_in[63]}),
		.sram(clk_mux_size3_95_sram[0:1]),
		.sram_inv(clk_mux_size3_95_sram_inv[0:1]),
		.out(chany_bottom_out[63]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_64 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[52:53]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[52:53]),
		.mem_out(clk_mux_size3_0_sram[0:1]),
		.mem_outb(clk_mux_size3_0_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_66 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[54:55]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[54:55]),
		.mem_out(clk_mux_size3_1_sram[0:1]),
		.mem_outb(clk_mux_size3_1_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_68 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[56:57]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[56:57]),
		.mem_out(clk_mux_size3_2_sram[0:1]),
		.mem_outb(clk_mux_size3_2_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_70 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[58:59]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[58:59]),
		.mem_out(clk_mux_size3_3_sram[0:1]),
		.mem_outb(clk_mux_size3_3_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_72 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[60:61]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[60:61]),
		.mem_out(clk_mux_size3_4_sram[0:1]),
		.mem_outb(clk_mux_size3_4_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_74 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[62:63]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[62:63]),
		.mem_out(clk_mux_size3_5_sram[0:1]),
		.mem_outb(clk_mux_size3_5_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_76 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[64:65]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[64:65]),
		.mem_out(clk_mux_size3_6_sram[0:1]),
		.mem_outb(clk_mux_size3_6_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_78 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[66:67]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[66:67]),
		.mem_out(clk_mux_size3_7_sram[0:1]),
		.mem_outb(clk_mux_size3_7_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_80 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[68:69]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[68:69]),
		.mem_out(clk_mux_size3_8_sram[0:1]),
		.mem_outb(clk_mux_size3_8_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_82 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[70:71]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[70:71]),
		.mem_out(clk_mux_size3_9_sram[0:1]),
		.mem_outb(clk_mux_size3_9_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_84 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[72:73]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[72:73]),
		.mem_out(clk_mux_size3_10_sram[0:1]),
		.mem_outb(clk_mux_size3_10_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_86 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[74:75]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[74:75]),
		.mem_out(clk_mux_size3_11_sram[0:1]),
		.mem_outb(clk_mux_size3_11_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_88 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[76:77]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[76:77]),
		.mem_out(clk_mux_size3_12_sram[0:1]),
		.mem_outb(clk_mux_size3_12_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_90 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[78:79]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[78:79]),
		.mem_out(clk_mux_size3_13_sram[0:1]),
		.mem_outb(clk_mux_size3_13_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_92 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[80:81]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[80:81]),
		.mem_out(clk_mux_size3_14_sram[0:1]),
		.mem_outb(clk_mux_size3_14_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_94 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[82:83]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[82:83]),
		.mem_out(clk_mux_size3_15_sram[0:1]),
		.mem_outb(clk_mux_size3_15_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_96 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[84:85]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[84:85]),
		.mem_out(clk_mux_size3_16_sram[0:1]),
		.mem_outb(clk_mux_size3_16_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_98 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[86:87]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[86:87]),
		.mem_out(clk_mux_size3_17_sram[0:1]),
		.mem_outb(clk_mux_size3_17_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_100 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[88:89]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[88:89]),
		.mem_out(clk_mux_size3_18_sram[0:1]),
		.mem_outb(clk_mux_size3_18_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_102 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[90:91]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[90:91]),
		.mem_out(clk_mux_size3_19_sram[0:1]),
		.mem_outb(clk_mux_size3_19_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_104 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[92:93]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[92:93]),
		.mem_out(clk_mux_size3_20_sram[0:1]),
		.mem_outb(clk_mux_size3_20_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_106 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[94:95]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[94:95]),
		.mem_out(clk_mux_size3_21_sram[0:1]),
		.mem_outb(clk_mux_size3_21_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_108 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[96:97]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[96:97]),
		.mem_out(clk_mux_size3_22_sram[0:1]),
		.mem_outb(clk_mux_size3_22_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_110 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[98:99]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[98:99]),
		.mem_out(clk_mux_size3_23_sram[0:1]),
		.mem_outb(clk_mux_size3_23_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_112 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[100:101]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[100:101]),
		.mem_out(clk_mux_size3_24_sram[0:1]),
		.mem_outb(clk_mux_size3_24_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_114 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[102:103]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[102:103]),
		.mem_out(clk_mux_size3_25_sram[0:1]),
		.mem_outb(clk_mux_size3_25_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_116 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[104:105]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[104:105]),
		.mem_out(clk_mux_size3_26_sram[0:1]),
		.mem_outb(clk_mux_size3_26_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_118 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[106:107]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[106:107]),
		.mem_out(clk_mux_size3_27_sram[0:1]),
		.mem_outb(clk_mux_size3_27_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_120 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[108:109]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[108:109]),
		.mem_out(clk_mux_size3_28_sram[0:1]),
		.mem_outb(clk_mux_size3_28_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_122 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[110:111]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[110:111]),
		.mem_out(clk_mux_size3_29_sram[0:1]),
		.mem_outb(clk_mux_size3_29_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_124 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[112:113]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[112:113]),
		.mem_out(clk_mux_size3_30_sram[0:1]),
		.mem_outb(clk_mux_size3_30_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_126 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[114:115]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[114:115]),
		.mem_out(clk_mux_size3_31_sram[0:1]),
		.mem_outb(clk_mux_size3_31_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_64 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[172:173]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[172:173]),
		.mem_out(clk_mux_size3_32_sram[0:1]),
		.mem_outb(clk_mux_size3_32_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_66 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[174:175]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[174:175]),
		.mem_out(clk_mux_size3_33_sram[0:1]),
		.mem_outb(clk_mux_size3_33_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_68 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[176:177]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[176:177]),
		.mem_out(clk_mux_size3_34_sram[0:1]),
		.mem_outb(clk_mux_size3_34_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_70 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[178:179]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[178:179]),
		.mem_out(clk_mux_size3_35_sram[0:1]),
		.mem_outb(clk_mux_size3_35_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_72 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[180:181]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[180:181]),
		.mem_out(clk_mux_size3_36_sram[0:1]),
		.mem_outb(clk_mux_size3_36_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_74 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[182:183]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[182:183]),
		.mem_out(clk_mux_size3_37_sram[0:1]),
		.mem_outb(clk_mux_size3_37_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_76 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[184:185]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[184:185]),
		.mem_out(clk_mux_size3_38_sram[0:1]),
		.mem_outb(clk_mux_size3_38_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_78 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[186:187]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[186:187]),
		.mem_out(clk_mux_size3_39_sram[0:1]),
		.mem_outb(clk_mux_size3_39_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_80 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[188:189]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[188:189]),
		.mem_out(clk_mux_size3_40_sram[0:1]),
		.mem_outb(clk_mux_size3_40_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_82 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[190:191]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[190:191]),
		.mem_out(clk_mux_size3_41_sram[0:1]),
		.mem_outb(clk_mux_size3_41_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_84 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[192:193]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[192:193]),
		.mem_out(clk_mux_size3_42_sram[0:1]),
		.mem_outb(clk_mux_size3_42_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_86 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[194:195]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[194:195]),
		.mem_out(clk_mux_size3_43_sram[0:1]),
		.mem_outb(clk_mux_size3_43_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_88 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[196:197]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[196:197]),
		.mem_out(clk_mux_size3_44_sram[0:1]),
		.mem_outb(clk_mux_size3_44_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_90 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[198:199]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[198:199]),
		.mem_out(clk_mux_size3_45_sram[0:1]),
		.mem_outb(clk_mux_size3_45_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_92 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[200:201]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[200:201]),
		.mem_out(clk_mux_size3_46_sram[0:1]),
		.mem_outb(clk_mux_size3_46_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_94 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[202:203]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[202:203]),
		.mem_out(clk_mux_size3_47_sram[0:1]),
		.mem_outb(clk_mux_size3_47_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_96 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[204:205]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[204:205]),
		.mem_out(clk_mux_size3_48_sram[0:1]),
		.mem_outb(clk_mux_size3_48_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_98 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[206:207]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[206:207]),
		.mem_out(clk_mux_size3_49_sram[0:1]),
		.mem_outb(clk_mux_size3_49_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_100 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[208:209]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[208:209]),
		.mem_out(clk_mux_size3_50_sram[0:1]),
		.mem_outb(clk_mux_size3_50_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_102 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[210:211]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[210:211]),
		.mem_out(clk_mux_size3_51_sram[0:1]),
		.mem_outb(clk_mux_size3_51_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_104 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[212:213]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[212:213]),
		.mem_out(clk_mux_size3_52_sram[0:1]),
		.mem_outb(clk_mux_size3_52_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_106 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[214:215]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[214:215]),
		.mem_out(clk_mux_size3_53_sram[0:1]),
		.mem_outb(clk_mux_size3_53_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_108 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[216:217]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[216:217]),
		.mem_out(clk_mux_size3_54_sram[0:1]),
		.mem_outb(clk_mux_size3_54_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_110 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[218:219]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[218:219]),
		.mem_out(clk_mux_size3_55_sram[0:1]),
		.mem_outb(clk_mux_size3_55_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_112 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[220:221]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[220:221]),
		.mem_out(clk_mux_size3_56_sram[0:1]),
		.mem_outb(clk_mux_size3_56_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_114 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[222:223]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[222:223]),
		.mem_out(clk_mux_size3_57_sram[0:1]),
		.mem_outb(clk_mux_size3_57_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_116 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[224:225]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[224:225]),
		.mem_out(clk_mux_size3_58_sram[0:1]),
		.mem_outb(clk_mux_size3_58_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_118 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[226:227]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[226:227]),
		.mem_out(clk_mux_size3_59_sram[0:1]),
		.mem_outb(clk_mux_size3_59_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_120 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[228:229]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[228:229]),
		.mem_out(clk_mux_size3_60_sram[0:1]),
		.mem_outb(clk_mux_size3_60_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_122 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[230:231]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[230:231]),
		.mem_out(clk_mux_size3_61_sram[0:1]),
		.mem_outb(clk_mux_size3_61_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_124 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[232:233]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[232:233]),
		.mem_out(clk_mux_size3_62_sram[0:1]),
		.mem_outb(clk_mux_size3_62_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_right_track_126 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[234:235]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[234:235]),
		.mem_out(clk_mux_size3_63_sram[0:1]),
		.mem_outb(clk_mux_size3_63_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_65 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[288:289]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[288:289]),
		.mem_out(clk_mux_size3_64_sram[0:1]),
		.mem_outb(clk_mux_size3_64_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_67 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[290:291]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[290:291]),
		.mem_out(clk_mux_size3_65_sram[0:1]),
		.mem_outb(clk_mux_size3_65_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_69 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[292:293]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[292:293]),
		.mem_out(clk_mux_size3_66_sram[0:1]),
		.mem_outb(clk_mux_size3_66_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_71 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[294:295]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[294:295]),
		.mem_out(clk_mux_size3_67_sram[0:1]),
		.mem_outb(clk_mux_size3_67_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_73 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[296:297]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[296:297]),
		.mem_out(clk_mux_size3_68_sram[0:1]),
		.mem_outb(clk_mux_size3_68_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_75 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[298:299]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[298:299]),
		.mem_out(clk_mux_size3_69_sram[0:1]),
		.mem_outb(clk_mux_size3_69_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_77 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[300:301]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[300:301]),
		.mem_out(clk_mux_size3_70_sram[0:1]),
		.mem_outb(clk_mux_size3_70_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_79 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[302:303]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[302:303]),
		.mem_out(clk_mux_size3_71_sram[0:1]),
		.mem_outb(clk_mux_size3_71_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_81 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[304:305]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[304:305]),
		.mem_out(clk_mux_size3_72_sram[0:1]),
		.mem_outb(clk_mux_size3_72_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_83 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[306:307]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[306:307]),
		.mem_out(clk_mux_size3_73_sram[0:1]),
		.mem_outb(clk_mux_size3_73_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_85 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[308:309]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[308:309]),
		.mem_out(clk_mux_size3_74_sram[0:1]),
		.mem_outb(clk_mux_size3_74_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_87 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[310:311]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[310:311]),
		.mem_out(clk_mux_size3_75_sram[0:1]),
		.mem_outb(clk_mux_size3_75_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_89 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[312:313]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[312:313]),
		.mem_out(clk_mux_size3_76_sram[0:1]),
		.mem_outb(clk_mux_size3_76_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_91 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[314:315]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[314:315]),
		.mem_out(clk_mux_size3_77_sram[0:1]),
		.mem_outb(clk_mux_size3_77_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_93 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[316:317]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[316:317]),
		.mem_out(clk_mux_size3_78_sram[0:1]),
		.mem_outb(clk_mux_size3_78_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_95 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[318:319]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[318:319]),
		.mem_out(clk_mux_size3_79_sram[0:1]),
		.mem_outb(clk_mux_size3_79_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_97 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[320:321]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[320:321]),
		.mem_out(clk_mux_size3_80_sram[0:1]),
		.mem_outb(clk_mux_size3_80_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_99 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[322:323]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[322:323]),
		.mem_out(clk_mux_size3_81_sram[0:1]),
		.mem_outb(clk_mux_size3_81_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_101 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[324:325]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[324:325]),
		.mem_out(clk_mux_size3_82_sram[0:1]),
		.mem_outb(clk_mux_size3_82_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_103 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[326:327]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[326:327]),
		.mem_out(clk_mux_size3_83_sram[0:1]),
		.mem_outb(clk_mux_size3_83_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_105 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[328:329]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[328:329]),
		.mem_out(clk_mux_size3_84_sram[0:1]),
		.mem_outb(clk_mux_size3_84_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_107 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[330:331]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[330:331]),
		.mem_out(clk_mux_size3_85_sram[0:1]),
		.mem_outb(clk_mux_size3_85_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_109 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[332:333]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[332:333]),
		.mem_out(clk_mux_size3_86_sram[0:1]),
		.mem_outb(clk_mux_size3_86_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_111 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[334:335]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[334:335]),
		.mem_out(clk_mux_size3_87_sram[0:1]),
		.mem_outb(clk_mux_size3_87_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_113 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[336:337]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[336:337]),
		.mem_out(clk_mux_size3_88_sram[0:1]),
		.mem_outb(clk_mux_size3_88_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_115 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[338:339]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[338:339]),
		.mem_out(clk_mux_size3_89_sram[0:1]),
		.mem_outb(clk_mux_size3_89_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_117 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[340:341]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[340:341]),
		.mem_out(clk_mux_size3_90_sram[0:1]),
		.mem_outb(clk_mux_size3_90_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_119 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[342:343]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[342:343]),
		.mem_out(clk_mux_size3_91_sram[0:1]),
		.mem_outb(clk_mux_size3_91_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_121 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[344:345]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[344:345]),
		.mem_out(clk_mux_size3_92_sram[0:1]),
		.mem_outb(clk_mux_size3_92_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_123 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[346:347]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[346:347]),
		.mem_out(clk_mux_size3_93_sram[0:1]),
		.mem_outb(clk_mux_size3_93_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_125 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[348:349]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[348:349]),
		.mem_out(clk_mux_size3_94_sram[0:1]),
		.mem_outb(clk_mux_size3_94_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_127 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[350:351]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[350:351]),
		.mem_out(clk_mux_size3_95_sram[0:1]),
		.mem_outb(clk_mux_size3_95_sram_inv[0:1]));

	sb_mux_size10 mux_right_track_0 (
		.in({chany_top_in[6], chany_top_in[26], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_, chany_bottom_in[6], chany_bottom_in[26:27], chanx_left_in[0]}),
		.sram(sb_mux_size10_0_sram[0:3]),
		.sram_inv(sb_mux_size10_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	sb_mux_size10 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[8], chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_, chany_bottom_in[8], chany_bottom_in[23], chany_bottom_in[28], chanx_left_in[1]}),
		.sram(sb_mux_size10_1_sram[0:3]),
		.sram_inv(sb_mux_size10_1_sram_inv[0:3]),
		.out(chanx_right_out[1]));

	sb_mux_size10 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[10], chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_, chany_bottom_in[10], chany_bottom_in[19], chany_bottom_in[29], chanx_left_in[2]}),
		.sram(sb_mux_size10_2_sram[0:3]),
		.sram_inv(sb_mux_size10_2_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	sb_mux_size10 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[12], chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_, chany_bottom_in[12], chany_bottom_in[15], chany_bottom_in[30], chanx_left_in[3]}),
		.sram(sb_mux_size10_3_sram[0:3]),
		.sram_inv(sb_mux_size10_3_sram_inv[0:3]),
		.out(chanx_right_out[3]));

	sb_mux_size10 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[6], chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_, chanx_right_in[0], chany_bottom_in[6], chany_bottom_in[26], chany_bottom_in[31]}),
		.sram(sb_mux_size10_4_sram[0:3]),
		.sram_inv(sb_mux_size10_4_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	sb_mux_size10 mux_left_track_3 (
		.in({chany_top_in[8], chany_top_in[28], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_, chanx_right_in[1], chany_bottom_in[0], chany_bottom_in[8], chany_bottom_in[28]}),
		.sram(sb_mux_size10_5_sram[0:3]),
		.sram_inv(sb_mux_size10_5_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	sb_mux_size10 mux_left_track_5 (
		.in({chany_top_in[10], chany_top_in[27], chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_, chanx_right_in[2], chany_bottom_in[1], chany_bottom_in[10], chany_bottom_in[29]}),
		.sram(sb_mux_size10_6_sram[0:3]),
		.sram_inv(sb_mux_size10_6_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	sb_mux_size10 mux_left_track_7 (
		.in({chany_top_in[12], chany_top_in[23], chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_, chanx_right_in[3], chany_bottom_in[2], chany_bottom_in[12], chany_bottom_in[30]}),
		.sram(sb_mux_size10_7_sram[0:3]),
		.sram_inv(sb_mux_size10_7_sram_inv[0:3]),
		.out(chanx_left_out[3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_right_track_0 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[116:119]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[116:119]),
		.mem_out(sb_mux_size10_0_sram[0:3]),
		.mem_outb(sb_mux_size10_0_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_right_track_2 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[120:123]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[120:123]),
		.mem_out(sb_mux_size10_1_sram[0:3]),
		.mem_outb(sb_mux_size10_1_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_right_track_4 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[124:127]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[124:127]),
		.mem_out(sb_mux_size10_2_sram[0:3]),
		.mem_outb(sb_mux_size10_2_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_right_track_6 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[128:131]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[128:131]),
		.mem_out(sb_mux_size10_3_sram[0:3]),
		.mem_outb(sb_mux_size10_3_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_left_track_1 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[352:355]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[352:355]),
		.mem_out(sb_mux_size10_4_sram[0:3]),
		.mem_outb(sb_mux_size10_4_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_left_track_3 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[356:359]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[356:359]),
		.mem_out(sb_mux_size10_5_sram[0:3]),
		.mem_outb(sb_mux_size10_5_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_left_track_5 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[360:363]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[360:363]),
		.mem_out(sb_mux_size10_6_sram[0:3]),
		.mem_outb(sb_mux_size10_6_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_left_track_7 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[364:367]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[364:367]),
		.mem_out(sb_mux_size10_7_sram[0:3]),
		.mem_outb(sb_mux_size10_7_sram_inv[0:3]));

	sb_mux_size8 mux_right_track_8 (
		.in({chany_top_in[3], chany_top_in[13], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_, chany_bottom_in[11], chany_bottom_in[13], chanx_left_in[4]}),
		.sram(sb_mux_size8_0_sram[0:3]),
		.sram_inv(sb_mux_size8_0_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	sb_mux_size8 mux_right_track_10 (
		.in({chany_top_in[4], chany_top_in[14], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_, chany_bottom_in[9], chany_bottom_in[14], chanx_left_in[5]}),
		.sram(sb_mux_size8_1_sram[0:3]),
		.sram_inv(sb_mux_size8_1_sram_inv[0:3]),
		.out(chanx_right_out[5]));

	sb_mux_size8 mux_right_track_48 (
		.in({chany_top_in[23:24], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_, chany_bottom_in[0], chany_bottom_in[24], chanx_left_in[27]}),
		.sram(sb_mux_size8_2_sram[0:3]),
		.sram_inv(sb_mux_size8_2_sram_inv[0:3]),
		.out(chanx_right_out[24]));

	sb_mux_size8 mux_right_track_56 (
		.in({chany_top_in[25], chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_, chany_bottom_in[25], chany_bottom_in[31], chanx_left_in[31]}),
		.sram(sb_mux_size8_3_sram[0:3]),
		.sram_inv(sb_mux_size8_3_sram_inv[0:3]),
		.out(chanx_right_out[28]));

	sb_mux_size8 mux_left_track_9 (
		.in({chany_top_in[13], chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_, chanx_right_in[4], chany_bottom_in[3], chany_bottom_in[13]}),
		.sram(sb_mux_size8_4_sram[0:3]),
		.sram_inv(sb_mux_size8_4_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	sb_mux_size8 mux_left_track_11 (
		.in({chany_top_in[14:15], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_, chanx_right_in[5], chany_bottom_in[4], chany_bottom_in[14]}),
		.sram(sb_mux_size8_5_sram[0:3]),
		.sram_inv(sb_mux_size8_5_sram_inv[0:3]),
		.out(chanx_left_out[5]));

	sb_mux_size8 mux_left_track_49 (
		.in({chany_top_in[2], chany_top_in[24], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_, chanx_right_in[27], chany_bottom_in[23:24]}),
		.sram(sb_mux_size8_6_sram[0:3]),
		.sram_inv(sb_mux_size8_6_sram_inv[0:3]),
		.out(chanx_left_out[24]));

	sb_mux_size8 mux_left_track_57 (
		.in({chany_top_in[1], chany_top_in[25], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_, chanx_right_in[31], chany_bottom_in[25], chany_bottom_in[27]}),
		.sram(sb_mux_size8_7_sram[0:3]),
		.sram_inv(sb_mux_size8_7_sram_inv[0:3]),
		.out(chanx_left_out[28]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_right_track_8 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[132:135]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[132:135]),
		.mem_out(sb_mux_size8_0_sram[0:3]),
		.mem_outb(sb_mux_size8_0_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_right_track_10 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[136:139]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[136:139]),
		.mem_out(sb_mux_size8_1_sram[0:3]),
		.mem_outb(sb_mux_size8_1_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_right_track_48 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[164:167]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[164:167]),
		.mem_out(sb_mux_size8_2_sram[0:3]),
		.mem_outb(sb_mux_size8_2_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_right_track_56 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[168:171]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[168:171]),
		.mem_out(sb_mux_size8_3_sram[0:3]),
		.mem_outb(sb_mux_size8_3_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_9 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[368:371]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[368:371]),
		.mem_out(sb_mux_size8_4_sram[0:3]),
		.mem_outb(sb_mux_size8_4_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_11 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[372:375]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[372:375]),
		.mem_out(sb_mux_size8_5_sram[0:3]),
		.mem_outb(sb_mux_size8_5_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_49 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[400:403]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[400:403]),
		.mem_out(sb_mux_size8_6_sram[0:3]),
		.mem_outb(sb_mux_size8_6_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_57 (
		.feedthrough_mem_in(sb_2__config_group_mem_size408_0_mem_out[404:407]),
		.feedthrough_mem_inb(sb_2__config_group_mem_size408_0_mem_outb[404:407]),
		.mem_out(sb_mux_size8_7_sram[0:3]),
		.mem_outb(sb_mux_size8_7_sram_inv[0:3]));

	sb_2__config_group_mem_size408 sb_2__config_group_mem_size408 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.mem_out(sb_2__config_group_mem_size408_0_mem_out[0:407]),
		.mem_outb(sb_2__config_group_mem_size408_0_mem_outb[0:407]),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for sb_2_ -----



