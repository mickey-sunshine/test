//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][5]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for sb_9_ -----
module sb_9_(chany_bottom_in,
             chany_bottom_out);
//----- INPUT PORTS -----
input [0:63] chany_bottom_in;
//----- OUTPUT PORTS -----
output [0:63] chany_bottom_out;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_9_ -----



