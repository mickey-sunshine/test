//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Fabric Netlist Summary
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ------ Include defines: preproc flags -----
`include "fpga_defines.v"

// ------ Include user-defined netlists -----
`include "./custom_modules/efpga_circuits.v"
// ------ Include primitive module netlists -----
`include "sub_module/inv_buf_passgate.v"
`include "sub_module/arch_encoder.v"
`include "sub_module/local_encoder.v"
`include "sub_module/mux_primitives.v"
`include "sub_module/muxes.v"
`include "sub_module/luts.v"
`include "sub_module/wires.v"
`include "sub_module/memories.v"
`include "sub_module/shift_register_banks.v"

// ------ Include logic block netlists -----
`include "lb/logical_tile_ckbuf_mode_ckbuf_physical_mode__ckbuf_core.v"
`include "lb/logical_tile_ckbuf_mode_ckbuf_.v"
`include "lb/logical_tile_clb_mode_clb_default_mode__fle_mode_fle_physical_mode__fabric_mode_fabric_default_mode___phy_fpga_adder_core.v"
`include "lb/logical_tile_clb_mode_clb_default_mode__fle_mode_fle_physical_mode__fabric_mode_fabric_default_mode__frac_logic_mode_frac_logic_default_mode__frac_lut5_arith_frac_lut5_arith.v"
`include "lb/logical_tile_clb_mode_clb_default_mode__fle_mode_fle_physical_mode__fabric_mode_fabric_default_mode__frac_logic.v"
`include "lb/logical_tile_clb_mode_clb_default_mode__fle_mode_fle_physical_mode__fabric_mode_fabric_default_mode__p_ff_p_ff.v"
`include "lb/logical_tile_clb_mode_clb_default_mode__fle_mode_fle_physical_mode__fabric.v"
`include "lb/logical_tile_clb_mode_clb_default_mode__fle.v"
`include "lb/logical_tile_clb_mode_clb_.v"
`include "lb/logical_tile_io_pi_mode_io_pi_physical_mode__pi_pad_mode_pi_pad_default_mode__io_pi_io_pi.v"
`include "lb/logical_tile_io_pi_mode_io_pi_physical_mode__pi_pad_mode_pi_pad_default_mode__p_io_scffi_p_io_scffi.v"
`include "lb/logical_tile_io_pi_mode_io_pi_physical_mode__pi_pad.v"
`include "lb/logical_tile_io_pi_mode_io_pi_.v"
`include "lb/logical_tile_io_pi_pdc_ecb1_mode_io_pi_pdc_ecb1_physical_mode__pi_pdc_ecb1_pad_mode_pi_pdc_ecb1_pad_default_mode__io_pi_pdc_ecb1_io_pi_pdc_ecb1.v"
`include "lb/logical_tile_io_pi_pdc_ecb1_mode_io_pi_pdc_ecb1_physical_mode__pi_pdc_ecb1_pad_mode_pi_pdc_ecb1_pad_default_mode__p_io_pdc_ecb1_scffi_p_io_pdc_ecb1_scffi.v"
`include "lb/logical_tile_io_pi_pdc_ecb1_mode_io_pi_pdc_ecb1_physical_mode__pi_pdc_ecb1_pad.v"
`include "lb/logical_tile_io_pi_pdc_ecb1_mode_io_pi_pdc_ecb1_.v"
`include "lb/logical_tile_io_po_mode_io_po_physical_mode__po_pad_mode_po_pad_default_mode__io_po_core.v"
`include "lb/logical_tile_io_po_mode_io_po_physical_mode__po_pad_mode_po_pad_default_mode__p_io_scffo_p_io_scffo.v"
`include "lb/logical_tile_io_po_mode_io_po_physical_mode__po_pad.v"
`include "lb/logical_tile_io_po_mode_io_po_.v"
`include "lb/logical_tile_io_po_cko_mode_io_po_cko_physical_mode__po_cko_pad_mode_po_cko_pad_default_mode__io_po_cko_core.v"
`include "lb/logical_tile_io_po_cko_mode_io_po_cko_physical_mode__po_cko_pad_mode_po_cko_pad_default_mode__p_io_cko_scffo_p_io_cko_scffo.v"
`include "lb/logical_tile_io_po_cko_mode_io_po_cko_physical_mode__po_cko_pad.v"
`include "lb/logical_tile_io_po_cko_mode_io_po_cko_.v"
`include "lb/logical_tile_pcnt_mode_pcnt_physical_mode___pcnt__pcnt.v"
`include "lb/logical_tile_pcnt_mode_pcnt_.v"
`include "lb/grid_clb.v"
`include "lb/grid_io_bottomL_bottom.v"
`include "lb/grid_io_leftL_left.v"
`include "lb/grid_io_rightL_right.v"
`include "lb/grid_io_topL_top.v"

// ------ Include routing module netlists -----
`include "routing/sb_0_.v"
`include "routing/sb_1_.v"
`include "routing/sb_2_.v"
`include "routing/sb_3_.v"
`include "routing/sb_4_.v"
`include "routing/sb_5_.v"
`include "routing/sb_6_.v"
`include "routing/sb_7_.v"
`include "routing/sb_8_.v"
`include "routing/sb_9_.v"
`include "routing/sb_10_.v"
`include "routing/sb_11_.v"
`include "routing/sb_12_.v"
`include "routing/sb_13_.v"
`include "routing/sb_14_.v"
`include "routing/cbx_0_.v"
`include "routing/cbx_1_.v"
`include "routing/cbx_2_.v"
`include "routing/cbx_3_.v"
`include "routing/cbx_4_.v"
`include "routing/cbx_5_.v"
`include "routing/cbx_6_.v"
`include "routing/cby_0_.v"
`include "routing/cby_1_.v"
`include "routing/cby_2_.v"
`include "routing/cby_3_.v"
`include "routing/cby_4_.v"
`include "routing/cby_5_.v"
`include "routing/cby_6_.v"

// ------ Include tile module netlists -----
`include "tile/tile_0__EMPTY_id7_.v"
`include "tile/tile_1__io_leftL_left_id8_.v"
`include "tile/tile_2__io_leftL_left_id9_.v"
`include "tile/tile_3__io_leftL_left_id10_.v"
`include "tile/tile_4__io_leftL_left_id11_.v"
`include "tile/tile_5__EMPTY_id0_.v"
`include "tile/tile_6__io_bottomL_bottom_id6_.v"
`include "tile/tile_7__clb_id12_.v"
`include "tile/tile_8__clb_id13_.v"
`include "tile/tile_9__io_topL_top_id1_.v"
`include "tile/tile_10__io_bottomL_bottom_id5_.v"
`include "tile/tile_11__clb_id14_.v"
`include "tile/tile_12__clb_id15_.v"
`include "tile/tile_13__EMPTY_id4_.v"
`include "tile/tile_14__io_rightL_right_id3_.v"
`include "tile/tile_15__io_rightL_right_id2_.v"

// ------ Include fabric top-level netlists -----
`include "fpga_core.v"
`include "fpga_top.v"

