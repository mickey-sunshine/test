//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for sb_6_ -----
module sb_6_(config_enable,
             prog_reset,
             prog_clk,
             chany_top_in,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_,
             top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_,
             top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_,
             top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_,
             top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_,
             chanx_right_in,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
             chany_bottom_in,
             chanx_left_in,
             left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
             left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
             left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
             left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
             left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
             left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
             left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
             left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
             ccff_head,
             chany_top_out,
             chanx_right_out,
             chany_bottom_out,
             chanx_left_out,
             ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:63] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_;
//----- INPUT PORTS -----
input [0:63] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:63] chany_bottom_in;
//----- INPUT PORTS -----
input [0:63] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:63] chany_top_out;
//----- OUTPUT PORTS -----
output [0:63] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:63] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:63] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] clk_mux_size3_0_sram;
wire [0:1] clk_mux_size3_0_sram_inv;
wire [0:1] clk_mux_size3_10_sram;
wire [0:1] clk_mux_size3_10_sram_inv;
wire [0:1] clk_mux_size3_11_sram;
wire [0:1] clk_mux_size3_11_sram_inv;
wire [0:1] clk_mux_size3_12_sram;
wire [0:1] clk_mux_size3_12_sram_inv;
wire [0:1] clk_mux_size3_13_sram;
wire [0:1] clk_mux_size3_13_sram_inv;
wire [0:1] clk_mux_size3_14_sram;
wire [0:1] clk_mux_size3_14_sram_inv;
wire [0:1] clk_mux_size3_15_sram;
wire [0:1] clk_mux_size3_15_sram_inv;
wire [0:1] clk_mux_size3_16_sram;
wire [0:1] clk_mux_size3_16_sram_inv;
wire [0:1] clk_mux_size3_17_sram;
wire [0:1] clk_mux_size3_17_sram_inv;
wire [0:1] clk_mux_size3_18_sram;
wire [0:1] clk_mux_size3_18_sram_inv;
wire [0:1] clk_mux_size3_19_sram;
wire [0:1] clk_mux_size3_19_sram_inv;
wire [0:1] clk_mux_size3_1_sram;
wire [0:1] clk_mux_size3_1_sram_inv;
wire [0:1] clk_mux_size3_20_sram;
wire [0:1] clk_mux_size3_20_sram_inv;
wire [0:1] clk_mux_size3_21_sram;
wire [0:1] clk_mux_size3_21_sram_inv;
wire [0:1] clk_mux_size3_22_sram;
wire [0:1] clk_mux_size3_22_sram_inv;
wire [0:1] clk_mux_size3_23_sram;
wire [0:1] clk_mux_size3_23_sram_inv;
wire [0:1] clk_mux_size3_24_sram;
wire [0:1] clk_mux_size3_24_sram_inv;
wire [0:1] clk_mux_size3_25_sram;
wire [0:1] clk_mux_size3_25_sram_inv;
wire [0:1] clk_mux_size3_26_sram;
wire [0:1] clk_mux_size3_26_sram_inv;
wire [0:1] clk_mux_size3_27_sram;
wire [0:1] clk_mux_size3_27_sram_inv;
wire [0:1] clk_mux_size3_28_sram;
wire [0:1] clk_mux_size3_28_sram_inv;
wire [0:1] clk_mux_size3_29_sram;
wire [0:1] clk_mux_size3_29_sram_inv;
wire [0:1] clk_mux_size3_2_sram;
wire [0:1] clk_mux_size3_2_sram_inv;
wire [0:1] clk_mux_size3_30_sram;
wire [0:1] clk_mux_size3_30_sram_inv;
wire [0:1] clk_mux_size3_31_sram;
wire [0:1] clk_mux_size3_31_sram_inv;
wire [0:1] clk_mux_size3_32_sram;
wire [0:1] clk_mux_size3_32_sram_inv;
wire [0:1] clk_mux_size3_33_sram;
wire [0:1] clk_mux_size3_33_sram_inv;
wire [0:1] clk_mux_size3_34_sram;
wire [0:1] clk_mux_size3_34_sram_inv;
wire [0:1] clk_mux_size3_35_sram;
wire [0:1] clk_mux_size3_35_sram_inv;
wire [0:1] clk_mux_size3_36_sram;
wire [0:1] clk_mux_size3_36_sram_inv;
wire [0:1] clk_mux_size3_37_sram;
wire [0:1] clk_mux_size3_37_sram_inv;
wire [0:1] clk_mux_size3_38_sram;
wire [0:1] clk_mux_size3_38_sram_inv;
wire [0:1] clk_mux_size3_39_sram;
wire [0:1] clk_mux_size3_39_sram_inv;
wire [0:1] clk_mux_size3_3_sram;
wire [0:1] clk_mux_size3_3_sram_inv;
wire [0:1] clk_mux_size3_40_sram;
wire [0:1] clk_mux_size3_40_sram_inv;
wire [0:1] clk_mux_size3_41_sram;
wire [0:1] clk_mux_size3_41_sram_inv;
wire [0:1] clk_mux_size3_42_sram;
wire [0:1] clk_mux_size3_42_sram_inv;
wire [0:1] clk_mux_size3_43_sram;
wire [0:1] clk_mux_size3_43_sram_inv;
wire [0:1] clk_mux_size3_44_sram;
wire [0:1] clk_mux_size3_44_sram_inv;
wire [0:1] clk_mux_size3_45_sram;
wire [0:1] clk_mux_size3_45_sram_inv;
wire [0:1] clk_mux_size3_46_sram;
wire [0:1] clk_mux_size3_46_sram_inv;
wire [0:1] clk_mux_size3_47_sram;
wire [0:1] clk_mux_size3_47_sram_inv;
wire [0:1] clk_mux_size3_48_sram;
wire [0:1] clk_mux_size3_48_sram_inv;
wire [0:1] clk_mux_size3_49_sram;
wire [0:1] clk_mux_size3_49_sram_inv;
wire [0:1] clk_mux_size3_4_sram;
wire [0:1] clk_mux_size3_4_sram_inv;
wire [0:1] clk_mux_size3_50_sram;
wire [0:1] clk_mux_size3_50_sram_inv;
wire [0:1] clk_mux_size3_51_sram;
wire [0:1] clk_mux_size3_51_sram_inv;
wire [0:1] clk_mux_size3_52_sram;
wire [0:1] clk_mux_size3_52_sram_inv;
wire [0:1] clk_mux_size3_53_sram;
wire [0:1] clk_mux_size3_53_sram_inv;
wire [0:1] clk_mux_size3_54_sram;
wire [0:1] clk_mux_size3_54_sram_inv;
wire [0:1] clk_mux_size3_55_sram;
wire [0:1] clk_mux_size3_55_sram_inv;
wire [0:1] clk_mux_size3_56_sram;
wire [0:1] clk_mux_size3_56_sram_inv;
wire [0:1] clk_mux_size3_57_sram;
wire [0:1] clk_mux_size3_57_sram_inv;
wire [0:1] clk_mux_size3_58_sram;
wire [0:1] clk_mux_size3_58_sram_inv;
wire [0:1] clk_mux_size3_59_sram;
wire [0:1] clk_mux_size3_59_sram_inv;
wire [0:1] clk_mux_size3_5_sram;
wire [0:1] clk_mux_size3_5_sram_inv;
wire [0:1] clk_mux_size3_60_sram;
wire [0:1] clk_mux_size3_60_sram_inv;
wire [0:1] clk_mux_size3_61_sram;
wire [0:1] clk_mux_size3_61_sram_inv;
wire [0:1] clk_mux_size3_62_sram;
wire [0:1] clk_mux_size3_62_sram_inv;
wire [0:1] clk_mux_size3_63_sram;
wire [0:1] clk_mux_size3_63_sram_inv;
wire [0:1] clk_mux_size3_6_sram;
wire [0:1] clk_mux_size3_6_sram_inv;
wire [0:1] clk_mux_size3_7_sram;
wire [0:1] clk_mux_size3_7_sram_inv;
wire [0:1] clk_mux_size3_8_sram;
wire [0:1] clk_mux_size3_8_sram_inv;
wire [0:1] clk_mux_size3_9_sram;
wire [0:1] clk_mux_size3_9_sram_inv;
wire [0:339] sb_6__config_group_mem_size340_0_mem_out;
wire [0:339] sb_6__config_group_mem_size340_0_mem_outb;
wire [0:3] sb_mux_size10_0_sram;
wire [0:3] sb_mux_size10_0_sram_inv;
wire [0:3] sb_mux_size10_10_sram;
wire [0:3] sb_mux_size10_10_sram_inv;
wire [0:3] sb_mux_size10_11_sram;
wire [0:3] sb_mux_size10_11_sram_inv;
wire [0:3] sb_mux_size10_1_sram;
wire [0:3] sb_mux_size10_1_sram_inv;
wire [0:3] sb_mux_size10_2_sram;
wire [0:3] sb_mux_size10_2_sram_inv;
wire [0:3] sb_mux_size10_3_sram;
wire [0:3] sb_mux_size10_3_sram_inv;
wire [0:3] sb_mux_size10_4_sram;
wire [0:3] sb_mux_size10_4_sram_inv;
wire [0:3] sb_mux_size10_5_sram;
wire [0:3] sb_mux_size10_5_sram_inv;
wire [0:3] sb_mux_size10_6_sram;
wire [0:3] sb_mux_size10_6_sram_inv;
wire [0:3] sb_mux_size10_7_sram;
wire [0:3] sb_mux_size10_7_sram_inv;
wire [0:3] sb_mux_size10_8_sram;
wire [0:3] sb_mux_size10_8_sram_inv;
wire [0:3] sb_mux_size10_9_sram;
wire [0:3] sb_mux_size10_9_sram_inv;
wire [0:3] sb_mux_size11_0_sram;
wire [0:3] sb_mux_size11_0_sram_inv;
wire [0:3] sb_mux_size11_1_sram;
wire [0:3] sb_mux_size11_1_sram_inv;
wire [0:3] sb_mux_size11_2_sram;
wire [0:3] sb_mux_size11_2_sram_inv;
wire [0:3] sb_mux_size11_3_sram;
wire [0:3] sb_mux_size11_3_sram_inv;
wire [0:3] sb_mux_size11_4_sram;
wire [0:3] sb_mux_size11_4_sram_inv;
wire [0:3] sb_mux_size11_5_sram;
wire [0:3] sb_mux_size11_5_sram_inv;
wire [0:3] sb_mux_size11_6_sram;
wire [0:3] sb_mux_size11_6_sram_inv;
wire [0:3] sb_mux_size11_7_sram;
wire [0:3] sb_mux_size11_7_sram_inv;
wire [0:2] sb_mux_size7_0_sram;
wire [0:2] sb_mux_size7_0_sram_inv;
wire [0:2] sb_mux_size7_10_sram;
wire [0:2] sb_mux_size7_10_sram_inv;
wire [0:2] sb_mux_size7_11_sram;
wire [0:2] sb_mux_size7_11_sram_inv;
wire [0:2] sb_mux_size7_1_sram;
wire [0:2] sb_mux_size7_1_sram_inv;
wire [0:2] sb_mux_size7_2_sram;
wire [0:2] sb_mux_size7_2_sram_inv;
wire [0:2] sb_mux_size7_3_sram;
wire [0:2] sb_mux_size7_3_sram_inv;
wire [0:2] sb_mux_size7_4_sram;
wire [0:2] sb_mux_size7_4_sram_inv;
wire [0:2] sb_mux_size7_5_sram;
wire [0:2] sb_mux_size7_5_sram_inv;
wire [0:2] sb_mux_size7_6_sram;
wire [0:2] sb_mux_size7_6_sram_inv;
wire [0:2] sb_mux_size7_7_sram;
wire [0:2] sb_mux_size7_7_sram_inv;
wire [0:2] sb_mux_size7_8_sram;
wire [0:2] sb_mux_size7_8_sram_inv;
wire [0:2] sb_mux_size7_9_sram;
wire [0:2] sb_mux_size7_9_sram_inv;
wire [0:3] sb_mux_size8_0_sram;
wire [0:3] sb_mux_size8_0_sram_inv;
wire [0:3] sb_mux_size8_1_sram;
wire [0:3] sb_mux_size8_1_sram_inv;
wire [0:3] sb_mux_size8_2_sram;
wire [0:3] sb_mux_size8_2_sram_inv;
wire [0:3] sb_mux_size8_3_sram;
wire [0:3] sb_mux_size8_3_sram_inv;
wire [0:3] sb_mux_size8_4_sram;
wire [0:3] sb_mux_size8_4_sram_inv;
wire [0:3] sb_mux_size8_5_sram;
wire [0:3] sb_mux_size8_5_sram_inv;
wire [0:3] sb_mux_size8_6_sram;
wire [0:3] sb_mux_size8_6_sram_inv;
wire [0:3] sb_mux_size8_7_sram;
wire [0:3] sb_mux_size8_7_sram_inv;
wire [0:3] sb_mux_size8_8_sram;
wire [0:3] sb_mux_size8_8_sram_inv;
wire [0:3] sb_mux_size8_9_sram;
wire [0:3] sb_mux_size8_9_sram_inv;
wire [0:3] sb_mux_size9_0_sram;
wire [0:3] sb_mux_size9_0_sram_inv;
wire [0:3] sb_mux_size9_10_sram;
wire [0:3] sb_mux_size9_10_sram_inv;
wire [0:3] sb_mux_size9_11_sram;
wire [0:3] sb_mux_size9_11_sram_inv;
wire [0:3] sb_mux_size9_12_sram;
wire [0:3] sb_mux_size9_12_sram_inv;
wire [0:3] sb_mux_size9_13_sram;
wire [0:3] sb_mux_size9_13_sram_inv;
wire [0:3] sb_mux_size9_1_sram;
wire [0:3] sb_mux_size9_1_sram_inv;
wire [0:3] sb_mux_size9_2_sram;
wire [0:3] sb_mux_size9_2_sram_inv;
wire [0:3] sb_mux_size9_3_sram;
wire [0:3] sb_mux_size9_3_sram_inv;
wire [0:3] sb_mux_size9_4_sram;
wire [0:3] sb_mux_size9_4_sram_inv;
wire [0:3] sb_mux_size9_5_sram;
wire [0:3] sb_mux_size9_5_sram_inv;
wire [0:3] sb_mux_size9_6_sram;
wire [0:3] sb_mux_size9_6_sram_inv;
wire [0:3] sb_mux_size9_7_sram;
wire [0:3] sb_mux_size9_7_sram_inv;
wire [0:3] sb_mux_size9_8_sram;
wire [0:3] sb_mux_size9_8_sram_inv;
wire [0:3] sb_mux_size9_9_sram;
wire [0:3] sb_mux_size9_9_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[32] = chanx_right_in[32];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[33];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[34];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[35];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[36] = chanx_right_in[36];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[37];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[38];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[39];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[40] = chanx_right_in[40];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[41];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[42];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[43];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[44] = chanx_right_in[44];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[45];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[46];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[47];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[48];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[49];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[50];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[51];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[52] = chanx_right_in[52];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[53];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[54];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[55];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[56] = chanx_right_in[56];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[57];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[58];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[59];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[60] = chanx_right_in[60];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[61];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[62];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[63];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[32] = chanx_left_in[32];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[33];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[34];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[35];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[36] = chanx_left_in[36];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[37];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[38];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[39];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[40] = chanx_left_in[40];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[41];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[42];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[43];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[44] = chanx_left_in[44];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[45];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[46];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[47];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[48] = chanx_left_in[48];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[49];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[50];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[51];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[52] = chanx_left_in[52];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[53];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[54];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[55];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[56] = chanx_left_in[56];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[57];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[58];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[59];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[60] = chanx_left_in[60];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[61];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[62];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[63];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size10 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chanx_right_in[1], chanx_right_in[6], chanx_right_in[26], chany_bottom_in[0], chanx_left_in[0], chanx_left_in[6], chanx_left_in[26]}),
		.sram(sb_mux_size10_0_sram[0:3]),
		.sram_inv(sb_mux_size10_0_sram_inv[0:3]),
		.out(chany_top_out[0]));

	sb_mux_size10 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chanx_right_in[2], chanx_right_in[8], chanx_right_in[28], chany_bottom_in[1], chanx_left_in[8], chanx_left_in[28], chanx_left_in[31]}),
		.sram(sb_mux_size10_1_sram[0:3]),
		.sram_inv(sb_mux_size10_1_sram_inv[0:3]),
		.out(chany_top_out[1]));

	sb_mux_size10 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chanx_right_in[3], chanx_right_in[10], chanx_right_in[29], chany_bottom_in[2], chanx_left_in[10], chanx_left_in[27], chanx_left_in[29]}),
		.sram(sb_mux_size10_2_sram[0:3]),
		.sram_inv(sb_mux_size10_2_sram_inv[0:3]),
		.out(chany_top_out[2]));

	sb_mux_size10 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chanx_right_in[9], chanx_right_in[16], chany_bottom_in[7], chanx_left_in[11], chanx_left_in[16]}),
		.sram(sb_mux_size10_3_sram[0:3]),
		.sram_inv(sb_mux_size10_3_sram_inv[0:3]),
		.out(chany_top_out[6]));

	sb_mux_size10 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chanx_right_in[11], chanx_right_in[17], chany_bottom_in[9], chanx_left_in[9], chanx_left_in[17]}),
		.sram(sb_mux_size10_4_sram[0:3]),
		.sram_inv(sb_mux_size10_4_sram_inv[0:3]),
		.out(chany_top_out[8]));

	sb_mux_size10 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chanx_right_in[15], chanx_right_in[18], chany_bottom_in[11], chanx_left_in[7], chanx_left_in[18]}),
		.sram(sb_mux_size10_5_sram[0:3]),
		.sram_inv(sb_mux_size10_5_sram_inv[0:3]),
		.out(chany_top_out[10]));

	sb_mux_size10 mux_bottom_track_1 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chany_top_in[0], chanx_right_in[6], chanx_right_in[26:27], chanx_left_in[1], chanx_left_in[6], chanx_left_in[26]}),
		.sram(sb_mux_size10_6_sram[0:3]),
		.sram_inv(sb_mux_size10_6_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	sb_mux_size10 mux_bottom_track_3 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chany_top_in[1], chanx_right_in[8], chanx_right_in[23], chanx_right_in[28], chanx_left_in[2], chanx_left_in[8], chanx_left_in[28]}),
		.sram(sb_mux_size10_7_sram[0:3]),
		.sram_inv(sb_mux_size10_7_sram_inv[0:3]),
		.out(chany_bottom_out[1]));

	sb_mux_size10 mux_bottom_track_5 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chany_top_in[2], chanx_right_in[10], chanx_right_in[19], chanx_right_in[29], chanx_left_in[3], chanx_left_in[10], chanx_left_in[29]}),
		.sram(sb_mux_size10_8_sram[0:3]),
		.sram_inv(sb_mux_size10_8_sram_inv[0:3]),
		.out(chany_bottom_out[2]));

	sb_mux_size10 mux_bottom_track_13 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chany_top_in[7], chanx_right_in[7], chanx_right_in[16], chanx_left_in[9], chanx_left_in[16]}),
		.sram(sb_mux_size10_9_sram[0:3]),
		.sram_inv(sb_mux_size10_9_sram_inv[0:3]),
		.out(chany_bottom_out[6]));

	sb_mux_size10 mux_bottom_track_17 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chany_top_in[9], chanx_right_in[5], chanx_right_in[17], chanx_left_in[11], chanx_left_in[17]}),
		.sram(sb_mux_size10_10_sram[0:3]),
		.sram_inv(sb_mux_size10_10_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	sb_mux_size10 mux_bottom_track_21 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chany_top_in[11], chanx_right_in[4], chanx_right_in[18], chanx_left_in[15], chanx_left_in[18]}),
		.sram(sb_mux_size10_11_sram[0:3]),
		.sram_inv(sb_mux_size10_11_sram_inv[0:3]),
		.out(chany_bottom_out[10]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_top_track_0 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[0:3]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[0:3]),
		.mem_out(sb_mux_size10_0_sram[0:3]),
		.mem_outb(sb_mux_size10_0_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_top_track_2 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[4:7]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[4:7]),
		.mem_out(sb_mux_size10_1_sram[0:3]),
		.mem_outb(sb_mux_size10_1_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_top_track_4 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[8:11]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[8:11]),
		.mem_out(sb_mux_size10_2_sram[0:3]),
		.mem_outb(sb_mux_size10_2_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_top_track_12 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[22:25]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[22:25]),
		.mem_out(sb_mux_size10_3_sram[0:3]),
		.mem_outb(sb_mux_size10_3_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_top_track_16 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[26:29]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[26:29]),
		.mem_out(sb_mux_size10_4_sram[0:3]),
		.mem_outb(sb_mux_size10_4_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_top_track_20 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[30:33]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[30:33]),
		.mem_out(sb_mux_size10_5_sram[0:3]),
		.mem_outb(sb_mux_size10_5_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_bottom_track_1 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[170:173]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[170:173]),
		.mem_out(sb_mux_size10_6_sram[0:3]),
		.mem_outb(sb_mux_size10_6_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_bottom_track_3 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[174:177]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[174:177]),
		.mem_out(sb_mux_size10_7_sram[0:3]),
		.mem_outb(sb_mux_size10_7_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_bottom_track_5 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[178:181]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[178:181]),
		.mem_out(sb_mux_size10_8_sram[0:3]),
		.mem_outb(sb_mux_size10_8_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_bottom_track_13 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[192:195]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[192:195]),
		.mem_out(sb_mux_size10_9_sram[0:3]),
		.mem_outb(sb_mux_size10_9_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_bottom_track_17 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[196:199]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[196:199]),
		.mem_out(sb_mux_size10_10_sram[0:3]),
		.mem_outb(sb_mux_size10_10_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_bottom_track_21 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[200:203]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[200:203]),
		.mem_out(sb_mux_size10_11_sram[0:3]),
		.mem_outb(sb_mux_size10_11_sram_inv[0:3]));

	sb_mux_size9 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_right_in[4], chanx_right_in[12], chanx_right_in[30], chany_bottom_in[3], chanx_left_in[12], chanx_left_in[23], chanx_left_in[30]}),
		.sram(sb_mux_size9_0_sram[0:3]),
		.sram_inv(sb_mux_size9_0_sram_inv[0:3]),
		.out(chany_top_out[3]));

	sb_mux_size9 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[10], chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, chany_bottom_in[10], chany_bottom_in[19], chany_bottom_in[29], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_left_in[2]}),
		.sram(sb_mux_size9_1_sram[0:3]),
		.sram_inv(sb_mux_size9_1_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	sb_mux_size9 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[12], chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_bottom_in[12], chany_bottom_in[15], chany_bottom_in[30], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_left_in[3]}),
		.sram(sb_mux_size9_2_sram[0:3]),
		.sram_inv(sb_mux_size9_2_sram_inv[0:3]),
		.out(chanx_right_out[3]));

	sb_mux_size9 mux_right_track_20 (
		.in({chany_top_in[9], chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[4], chany_bottom_in[18], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[11]}),
		.sram(sb_mux_size9_3_sram[0:3]),
		.sram_inv(sb_mux_size9_3_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	sb_mux_size9 mux_right_track_24 (
		.in({chany_top_in[11], chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[3], chany_bottom_in[20], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[15]}),
		.sram(sb_mux_size9_4_sram[0:3]),
		.sram_inv(sb_mux_size9_4_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	sb_mux_size9 mux_right_track_32 (
		.in({chany_top_in[15], chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[2], chany_bottom_in[21], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[19]}),
		.sram(sb_mux_size9_5_sram[0:3]),
		.sram_inv(sb_mux_size9_5_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	sb_mux_size9 mux_right_track_40 (
		.in({chany_top_in[19], chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[1], chany_bottom_in[22], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[23]}),
		.sram(sb_mux_size9_6_sram[0:3]),
		.sram_inv(sb_mux_size9_6_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	sb_mux_size9 mux_bottom_track_7 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chany_top_in[3], chanx_right_in[12], chanx_right_in[15], chanx_right_in[30], chanx_left_in[4], chanx_left_in[12], chanx_left_in[30]}),
		.sram(sb_mux_size9_7_sram[0:3]),
		.sram_inv(sb_mux_size9_7_sram_inv[0:3]),
		.out(chany_bottom_out[3]));

	sb_mux_size9 mux_left_track_5 (
		.in({chany_top_in[10], chany_top_in[27], chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_right_in[2], chany_bottom_in[1], chany_bottom_in[10], chany_bottom_in[29], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_}),
		.sram(sb_mux_size9_8_sram[0:3]),
		.sram_inv(sb_mux_size9_8_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	sb_mux_size9 mux_left_track_7 (
		.in({chany_top_in[12], chany_top_in[23], chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[3], chany_bottom_in[2], chany_bottom_in[12], chany_bottom_in[30], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_}),
		.sram(sb_mux_size9_9_sram[0:3]),
		.sram_inv(sb_mux_size9_9_sram_inv[0:3]),
		.out(chanx_left_out[3]));

	sb_mux_size9 mux_left_track_21 (
		.in({chany_top_in[7], chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[11], chany_bottom_in[9], chany_bottom_in[18], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(sb_mux_size9_10_sram[0:3]),
		.sram_inv(sb_mux_size9_10_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	sb_mux_size9 mux_left_track_25 (
		.in({chany_top_in[5], chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[15], chany_bottom_in[11], chany_bottom_in[20], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(sb_mux_size9_11_sram[0:3]),
		.sram_inv(sb_mux_size9_11_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	sb_mux_size9 mux_left_track_33 (
		.in({chany_top_in[4], chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[19], chany_bottom_in[15], chany_bottom_in[21], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_}),
		.sram(sb_mux_size9_12_sram[0:3]),
		.sram_inv(sb_mux_size9_12_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	sb_mux_size9 mux_left_track_41 (
		.in({chany_top_in[3], chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[23], chany_bottom_in[19], chany_bottom_in[22], left_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_}),
		.sram(sb_mux_size9_13_sram[0:3]),
		.sram_inv(sb_mux_size9_13_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_6 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[12:15]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[12:15]),
		.mem_out(sb_mux_size9_0_sram[0:3]),
		.mem_outb(sb_mux_size9_0_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_4 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[126:129]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[126:129]),
		.mem_out(sb_mux_size9_1_sram[0:3]),
		.mem_outb(sb_mux_size9_1_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_6 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[130:133]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[130:133]),
		.mem_out(sb_mux_size9_2_sram[0:3]),
		.mem_outb(sb_mux_size9_2_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_20 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[148:151]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[148:151]),
		.mem_out(sb_mux_size9_3_sram[0:3]),
		.mem_outb(sb_mux_size9_3_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_24 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[152:155]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[152:155]),
		.mem_out(sb_mux_size9_4_sram[0:3]),
		.mem_outb(sb_mux_size9_4_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_32 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[156:159]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[156:159]),
		.mem_out(sb_mux_size9_5_sram[0:3]),
		.mem_outb(sb_mux_size9_5_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_right_track_40 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[160:163]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[160:163]),
		.mem_out(sb_mux_size9_6_sram[0:3]),
		.mem_outb(sb_mux_size9_6_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_bottom_track_7 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[182:185]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[182:185]),
		.mem_out(sb_mux_size9_7_sram[0:3]),
		.mem_outb(sb_mux_size9_7_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_5 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[296:299]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[296:299]),
		.mem_out(sb_mux_size9_8_sram[0:3]),
		.mem_outb(sb_mux_size9_8_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_7 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[300:303]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[300:303]),
		.mem_out(sb_mux_size9_9_sram[0:3]),
		.mem_outb(sb_mux_size9_9_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_21 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[318:321]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[318:321]),
		.mem_out(sb_mux_size9_10_sram[0:3]),
		.mem_outb(sb_mux_size9_10_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_25 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[322:325]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[322:325]),
		.mem_out(sb_mux_size9_11_sram[0:3]),
		.mem_outb(sb_mux_size9_11_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_33 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[326:329]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[326:329]),
		.mem_out(sb_mux_size9_12_sram[0:3]),
		.mem_outb(sb_mux_size9_12_sram_inv[0:3]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_left_track_41 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[330:333]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[330:333]),
		.mem_out(sb_mux_size9_13_sram[0:3]),
		.mem_outb(sb_mux_size9_13_sram_inv[0:3]));

	sb_mux_size7 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_right_in[5], chanx_right_in[13], chany_bottom_in[4], chanx_left_in[13], chanx_left_in[19]}),
		.sram(sb_mux_size7_0_sram[0:2]),
		.sram_inv(sb_mux_size7_0_sram_inv[0:2]),
		.out(chany_top_out[4]));

	sb_mux_size7 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[7], chanx_right_in[14], chany_bottom_in[5], chanx_left_in[14:15]}),
		.sram(sb_mux_size7_1_sram[0:2]),
		.sram_inv(sb_mux_size7_1_sram_inv[0:2]),
		.out(chany_top_out[5]));

	sb_mux_size7 mux_right_track_8 (
		.in({chany_top_in[3], chany_top_in[13], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_bottom_in[11], chany_bottom_in[13], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_left_in[4]}),
		.sram(sb_mux_size7_2_sram[0:2]),
		.sram_inv(sb_mux_size7_2_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	sb_mux_size7 mux_right_track_10 (
		.in({chany_top_in[4], chany_top_in[14], right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chany_bottom_in[9], chany_bottom_in[14], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[5]}),
		.sram(sb_mux_size7_3_sram[0:2]),
		.sram_inv(sb_mux_size7_3_sram_inv[0:2]),
		.out(chanx_right_out[5]));

	sb_mux_size7 mux_right_track_48 (
		.in({chany_top_in[23:24], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chany_bottom_in[0], chany_bottom_in[24], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_left_in[27]}),
		.sram(sb_mux_size7_4_sram[0:2]),
		.sram_inv(sb_mux_size7_4_sram_inv[0:2]),
		.out(chanx_right_out[24]));

	sb_mux_size7 mux_right_track_56 (
		.in({chany_top_in[25], chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chany_bottom_in[25], chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_left_in[31]}),
		.sram(sb_mux_size7_5_sram[0:2]),
		.sram_inv(sb_mux_size7_5_sram_inv[0:2]),
		.out(chanx_right_out[28]));

	sb_mux_size7 mux_bottom_track_9 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chany_top_in[4], chanx_right_in[11], chanx_right_in[13], chanx_left_in[5], chanx_left_in[13]}),
		.sram(sb_mux_size7_6_sram[0:2]),
		.sram_inv(sb_mux_size7_6_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	sb_mux_size7 mux_bottom_track_11 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chany_top_in[5], chanx_right_in[9], chanx_right_in[14], chanx_left_in[7], chanx_left_in[14]}),
		.sram(sb_mux_size7_7_sram[0:2]),
		.sram_inv(sb_mux_size7_7_sram_inv[0:2]),
		.out(chany_bottom_out[5]));

	sb_mux_size7 mux_left_track_9 (
		.in({chany_top_in[13], chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[4], chany_bottom_in[3], chany_bottom_in[13], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(sb_mux_size7_8_sram[0:2]),
		.sram_inv(sb_mux_size7_8_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	sb_mux_size7 mux_left_track_11 (
		.in({chany_top_in[14:15], right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[5], chany_bottom_in[4], chany_bottom_in[14], left_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_}),
		.sram(sb_mux_size7_9_sram[0:2]),
		.sram_inv(sb_mux_size7_9_sram_inv[0:2]),
		.out(chanx_left_out[5]));

	sb_mux_size7 mux_left_track_49 (
		.in({chany_top_in[2], chany_top_in[24], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[27], chany_bottom_in[23:24], left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_}),
		.sram(sb_mux_size7_10_sram[0:2]),
		.sram_inv(sb_mux_size7_10_sram_inv[0:2]),
		.out(chanx_left_out[24]));

	sb_mux_size7 mux_left_track_57 (
		.in({chany_top_in[1], chany_top_in[25], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[31], chany_bottom_in[25], chany_bottom_in[27], left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_}),
		.sram(sb_mux_size7_11_sram[0:2]),
		.sram_inv(sb_mux_size7_11_sram_inv[0:2]),
		.out(chanx_left_out[28]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_8 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[16:18]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[16:18]),
		.mem_out(sb_mux_size7_0_sram[0:2]),
		.mem_outb(sb_mux_size7_0_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_10 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[19:21]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[19:21]),
		.mem_out(sb_mux_size7_1_sram[0:2]),
		.mem_outb(sb_mux_size7_1_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_right_track_8 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[134:136]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[134:136]),
		.mem_out(sb_mux_size7_2_sram[0:2]),
		.mem_outb(sb_mux_size7_2_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_right_track_10 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[137:139]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[137:139]),
		.mem_out(sb_mux_size7_3_sram[0:2]),
		.mem_outb(sb_mux_size7_3_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_right_track_48 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[164:166]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[164:166]),
		.mem_out(sb_mux_size7_4_sram[0:2]),
		.mem_outb(sb_mux_size7_4_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_right_track_56 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[167:169]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[167:169]),
		.mem_out(sb_mux_size7_5_sram[0:2]),
		.mem_outb(sb_mux_size7_5_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_9 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[186:188]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[186:188]),
		.mem_out(sb_mux_size7_6_sram[0:2]),
		.mem_outb(sb_mux_size7_6_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_11 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[189:191]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[189:191]),
		.mem_out(sb_mux_size7_7_sram[0:2]),
		.mem_outb(sb_mux_size7_7_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_9 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[304:306]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[304:306]),
		.mem_out(sb_mux_size7_8_sram[0:2]),
		.mem_outb(sb_mux_size7_8_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_11 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[307:309]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[307:309]),
		.mem_out(sb_mux_size7_9_sram[0:2]),
		.mem_outb(sb_mux_size7_9_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_49 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[334:336]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[334:336]),
		.mem_out(sb_mux_size7_10_sram[0:2]),
		.mem_outb(sb_mux_size7_10_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_57 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[337:339]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[337:339]),
		.mem_out(sb_mux_size7_11_sram[0:2]),
		.mem_outb(sb_mux_size7_11_sram_inv[0:2]));

	sb_mux_size8 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_right_in[19:20], chany_bottom_in[15], chanx_left_in[5], chanx_left_in[20]}),
		.sram(sb_mux_size8_0_sram[0:3]),
		.sram_inv(sb_mux_size8_0_sram_inv[0:3]),
		.out(chany_top_out[12]));

	sb_mux_size8 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_right_in[21], chanx_right_in[23], chany_bottom_in[19], chanx_left_in[4], chanx_left_in[21]}),
		.sram(sb_mux_size8_1_sram[0:3]),
		.sram_inv(sb_mux_size8_1_sram_inv[0:3]),
		.out(chany_top_out[16]));

	sb_mux_size8 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chanx_right_in[22], chanx_right_in[27], chany_bottom_in[23], chanx_left_in[3], chanx_left_in[22]}),
		.sram(sb_mux_size8_2_sram[0:3]),
		.sram_inv(sb_mux_size8_2_sram_inv[0:3]),
		.out(chany_top_out[20]));

	sb_mux_size8 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chanx_right_in[24], chanx_right_in[31], chany_bottom_in[27], chanx_left_in[2], chanx_left_in[24]}),
		.sram(sb_mux_size8_3_sram[0:3]),
		.sram_inv(sb_mux_size8_3_sram_inv[0:3]),
		.out(chany_top_out[24]));

	sb_mux_size8 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chanx_right_in[0], chanx_right_in[25], chany_bottom_in[31], chanx_left_in[1], chanx_left_in[25]}),
		.sram(sb_mux_size8_4_sram[0:3]),
		.sram_inv(sb_mux_size8_4_sram_inv[0:3]),
		.out(chany_top_out[28]));

	sb_mux_size8 mux_bottom_track_25 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chany_top_in[15], chanx_right_in[3], chanx_right_in[20], chanx_left_in[19:20]}),
		.sram(sb_mux_size8_5_sram[0:3]),
		.sram_inv(sb_mux_size8_5_sram_inv[0:3]),
		.out(chany_bottom_out[12]));

	sb_mux_size8 mux_bottom_track_33 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chany_top_in[19], chanx_right_in[2], chanx_right_in[21], chanx_left_in[21], chanx_left_in[23]}),
		.sram(sb_mux_size8_6_sram[0:3]),
		.sram_inv(sb_mux_size8_6_sram_inv[0:3]),
		.out(chany_bottom_out[16]));

	sb_mux_size8 mux_bottom_track_41 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chany_top_in[23], chanx_right_in[1], chanx_right_in[22], chanx_left_in[22], chanx_left_in[27]}),
		.sram(sb_mux_size8_7_sram[0:3]),
		.sram_inv(sb_mux_size8_7_sram_inv[0:3]),
		.out(chany_bottom_out[20]));

	sb_mux_size8 mux_bottom_track_49 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chany_top_in[27], chanx_right_in[0], chanx_right_in[24], chanx_left_in[24], chanx_left_in[31]}),
		.sram(sb_mux_size8_8_sram[0:3]),
		.sram_inv(sb_mux_size8_8_sram_inv[0:3]),
		.out(chany_bottom_out[24]));

	sb_mux_size8 mux_bottom_track_57 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chany_top_in[31], chanx_right_in[25], chanx_right_in[31], chanx_left_in[0], chanx_left_in[25]}),
		.sram(sb_mux_size8_9_sram[0:3]),
		.sram_inv(sb_mux_size8_9_sram_inv[0:3]),
		.out(chany_bottom_out[28]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_24 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[34:37]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[34:37]),
		.mem_out(sb_mux_size8_0_sram[0:3]),
		.mem_outb(sb_mux_size8_0_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_32 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[38:41]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[38:41]),
		.mem_out(sb_mux_size8_1_sram[0:3]),
		.mem_outb(sb_mux_size8_1_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_40 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[42:45]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[42:45]),
		.mem_out(sb_mux_size8_2_sram[0:3]),
		.mem_outb(sb_mux_size8_2_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_48 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[46:49]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[46:49]),
		.mem_out(sb_mux_size8_3_sram[0:3]),
		.mem_outb(sb_mux_size8_3_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_56 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[50:53]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[50:53]),
		.mem_out(sb_mux_size8_4_sram[0:3]),
		.mem_outb(sb_mux_size8_4_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_25 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[204:207]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[204:207]),
		.mem_out(sb_mux_size8_5_sram[0:3]),
		.mem_outb(sb_mux_size8_5_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_33 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[208:211]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[208:211]),
		.mem_out(sb_mux_size8_6_sram[0:3]),
		.mem_outb(sb_mux_size8_6_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_41 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[212:215]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[212:215]),
		.mem_out(sb_mux_size8_7_sram[0:3]),
		.mem_outb(sb_mux_size8_7_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_49 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[216:219]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[216:219]),
		.mem_out(sb_mux_size8_8_sram[0:3]),
		.mem_outb(sb_mux_size8_8_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_57 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[220:223]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[220:223]),
		.mem_out(sb_mux_size8_9_sram[0:3]),
		.mem_outb(sb_mux_size8_9_sram_inv[0:3]));

	clk_mux_size3 mux_top_track_64 (
		.in({chanx_right_in[32], chany_bottom_in[32], chanx_left_in[32]}),
		.sram(clk_mux_size3_0_sram[0:1]),
		.sram_inv(clk_mux_size3_0_sram_inv[0:1]),
		.out(chany_top_out[32]));

	clk_mux_size3 mux_top_track_66 (
		.in({chanx_right_in[33], chany_bottom_in[33], chanx_left_in[33]}),
		.sram(clk_mux_size3_1_sram[0:1]),
		.sram_inv(clk_mux_size3_1_sram_inv[0:1]),
		.out(chany_top_out[33]));

	clk_mux_size3 mux_top_track_68 (
		.in({chanx_right_in[34], chany_bottom_in[34], chanx_left_in[34]}),
		.sram(clk_mux_size3_2_sram[0:1]),
		.sram_inv(clk_mux_size3_2_sram_inv[0:1]),
		.out(chany_top_out[34]));

	clk_mux_size3 mux_top_track_70 (
		.in({chanx_right_in[35], chany_bottom_in[35], chanx_left_in[35]}),
		.sram(clk_mux_size3_3_sram[0:1]),
		.sram_inv(clk_mux_size3_3_sram_inv[0:1]),
		.out(chany_top_out[35]));

	clk_mux_size3 mux_top_track_72 (
		.in({chanx_right_in[36], chany_bottom_in[36], chanx_left_in[36]}),
		.sram(clk_mux_size3_4_sram[0:1]),
		.sram_inv(clk_mux_size3_4_sram_inv[0:1]),
		.out(chany_top_out[36]));

	clk_mux_size3 mux_top_track_74 (
		.in({chanx_right_in[37], chany_bottom_in[37], chanx_left_in[37]}),
		.sram(clk_mux_size3_5_sram[0:1]),
		.sram_inv(clk_mux_size3_5_sram_inv[0:1]),
		.out(chany_top_out[37]));

	clk_mux_size3 mux_top_track_76 (
		.in({chanx_right_in[38], chany_bottom_in[38], chanx_left_in[38]}),
		.sram(clk_mux_size3_6_sram[0:1]),
		.sram_inv(clk_mux_size3_6_sram_inv[0:1]),
		.out(chany_top_out[38]));

	clk_mux_size3 mux_top_track_78 (
		.in({chanx_right_in[39], chany_bottom_in[39], chanx_left_in[39]}),
		.sram(clk_mux_size3_7_sram[0:1]),
		.sram_inv(clk_mux_size3_7_sram_inv[0:1]),
		.out(chany_top_out[39]));

	clk_mux_size3 mux_top_track_80 (
		.in({chanx_right_in[40], chany_bottom_in[40], chanx_left_in[40]}),
		.sram(clk_mux_size3_8_sram[0:1]),
		.sram_inv(clk_mux_size3_8_sram_inv[0:1]),
		.out(chany_top_out[40]));

	clk_mux_size3 mux_top_track_82 (
		.in({chanx_right_in[41], chany_bottom_in[41], chanx_left_in[41]}),
		.sram(clk_mux_size3_9_sram[0:1]),
		.sram_inv(clk_mux_size3_9_sram_inv[0:1]),
		.out(chany_top_out[41]));

	clk_mux_size3 mux_top_track_84 (
		.in({chanx_right_in[42], chany_bottom_in[42], chanx_left_in[42]}),
		.sram(clk_mux_size3_10_sram[0:1]),
		.sram_inv(clk_mux_size3_10_sram_inv[0:1]),
		.out(chany_top_out[42]));

	clk_mux_size3 mux_top_track_86 (
		.in({chanx_right_in[43], chany_bottom_in[43], chanx_left_in[43]}),
		.sram(clk_mux_size3_11_sram[0:1]),
		.sram_inv(clk_mux_size3_11_sram_inv[0:1]),
		.out(chany_top_out[43]));

	clk_mux_size3 mux_top_track_88 (
		.in({chanx_right_in[44], chany_bottom_in[44], chanx_left_in[44]}),
		.sram(clk_mux_size3_12_sram[0:1]),
		.sram_inv(clk_mux_size3_12_sram_inv[0:1]),
		.out(chany_top_out[44]));

	clk_mux_size3 mux_top_track_90 (
		.in({chanx_right_in[45], chany_bottom_in[45], chanx_left_in[45]}),
		.sram(clk_mux_size3_13_sram[0:1]),
		.sram_inv(clk_mux_size3_13_sram_inv[0:1]),
		.out(chany_top_out[45]));

	clk_mux_size3 mux_top_track_92 (
		.in({chanx_right_in[46], chany_bottom_in[46], chanx_left_in[46]}),
		.sram(clk_mux_size3_14_sram[0:1]),
		.sram_inv(clk_mux_size3_14_sram_inv[0:1]),
		.out(chany_top_out[46]));

	clk_mux_size3 mux_top_track_94 (
		.in({chanx_right_in[47], chany_bottom_in[47], chanx_left_in[47]}),
		.sram(clk_mux_size3_15_sram[0:1]),
		.sram_inv(clk_mux_size3_15_sram_inv[0:1]),
		.out(chany_top_out[47]));

	clk_mux_size3 mux_top_track_96 (
		.in({chanx_right_in[48], chany_bottom_in[48], chanx_left_in[48]}),
		.sram(clk_mux_size3_16_sram[0:1]),
		.sram_inv(clk_mux_size3_16_sram_inv[0:1]),
		.out(chany_top_out[48]));

	clk_mux_size3 mux_top_track_98 (
		.in({chanx_right_in[49], chany_bottom_in[49], chanx_left_in[49]}),
		.sram(clk_mux_size3_17_sram[0:1]),
		.sram_inv(clk_mux_size3_17_sram_inv[0:1]),
		.out(chany_top_out[49]));

	clk_mux_size3 mux_top_track_100 (
		.in({chanx_right_in[50], chany_bottom_in[50], chanx_left_in[50]}),
		.sram(clk_mux_size3_18_sram[0:1]),
		.sram_inv(clk_mux_size3_18_sram_inv[0:1]),
		.out(chany_top_out[50]));

	clk_mux_size3 mux_top_track_102 (
		.in({chanx_right_in[51], chany_bottom_in[51], chanx_left_in[51]}),
		.sram(clk_mux_size3_19_sram[0:1]),
		.sram_inv(clk_mux_size3_19_sram_inv[0:1]),
		.out(chany_top_out[51]));

	clk_mux_size3 mux_top_track_104 (
		.in({chanx_right_in[52], chany_bottom_in[52], chanx_left_in[52]}),
		.sram(clk_mux_size3_20_sram[0:1]),
		.sram_inv(clk_mux_size3_20_sram_inv[0:1]),
		.out(chany_top_out[52]));

	clk_mux_size3 mux_top_track_106 (
		.in({chanx_right_in[53], chany_bottom_in[53], chanx_left_in[53]}),
		.sram(clk_mux_size3_21_sram[0:1]),
		.sram_inv(clk_mux_size3_21_sram_inv[0:1]),
		.out(chany_top_out[53]));

	clk_mux_size3 mux_top_track_108 (
		.in({chanx_right_in[54], chany_bottom_in[54], chanx_left_in[54]}),
		.sram(clk_mux_size3_22_sram[0:1]),
		.sram_inv(clk_mux_size3_22_sram_inv[0:1]),
		.out(chany_top_out[54]));

	clk_mux_size3 mux_top_track_110 (
		.in({chanx_right_in[55], chany_bottom_in[55], chanx_left_in[55]}),
		.sram(clk_mux_size3_23_sram[0:1]),
		.sram_inv(clk_mux_size3_23_sram_inv[0:1]),
		.out(chany_top_out[55]));

	clk_mux_size3 mux_top_track_112 (
		.in({chanx_right_in[56], chany_bottom_in[56], chanx_left_in[56]}),
		.sram(clk_mux_size3_24_sram[0:1]),
		.sram_inv(clk_mux_size3_24_sram_inv[0:1]),
		.out(chany_top_out[56]));

	clk_mux_size3 mux_top_track_114 (
		.in({chanx_right_in[57], chany_bottom_in[57], chanx_left_in[57]}),
		.sram(clk_mux_size3_25_sram[0:1]),
		.sram_inv(clk_mux_size3_25_sram_inv[0:1]),
		.out(chany_top_out[57]));

	clk_mux_size3 mux_top_track_116 (
		.in({chanx_right_in[58], chany_bottom_in[58], chanx_left_in[58]}),
		.sram(clk_mux_size3_26_sram[0:1]),
		.sram_inv(clk_mux_size3_26_sram_inv[0:1]),
		.out(chany_top_out[58]));

	clk_mux_size3 mux_top_track_118 (
		.in({chanx_right_in[59], chany_bottom_in[59], chanx_left_in[59]}),
		.sram(clk_mux_size3_27_sram[0:1]),
		.sram_inv(clk_mux_size3_27_sram_inv[0:1]),
		.out(chany_top_out[59]));

	clk_mux_size3 mux_top_track_120 (
		.in({chanx_right_in[60], chany_bottom_in[60], chanx_left_in[60]}),
		.sram(clk_mux_size3_28_sram[0:1]),
		.sram_inv(clk_mux_size3_28_sram_inv[0:1]),
		.out(chany_top_out[60]));

	clk_mux_size3 mux_top_track_122 (
		.in({chanx_right_in[61], chany_bottom_in[61], chanx_left_in[61]}),
		.sram(clk_mux_size3_29_sram[0:1]),
		.sram_inv(clk_mux_size3_29_sram_inv[0:1]),
		.out(chany_top_out[61]));

	clk_mux_size3 mux_top_track_124 (
		.in({chanx_right_in[62], chany_bottom_in[62], chanx_left_in[62]}),
		.sram(clk_mux_size3_30_sram[0:1]),
		.sram_inv(clk_mux_size3_30_sram_inv[0:1]),
		.out(chany_top_out[62]));

	clk_mux_size3 mux_top_track_126 (
		.in({chanx_right_in[63], chany_bottom_in[63], chanx_left_in[63]}),
		.sram(clk_mux_size3_31_sram[0:1]),
		.sram_inv(clk_mux_size3_31_sram_inv[0:1]),
		.out(chany_top_out[63]));

	clk_mux_size3 mux_bottom_track_65 (
		.in({chany_top_in[32], chanx_right_in[32], chanx_left_in[32]}),
		.sram(clk_mux_size3_32_sram[0:1]),
		.sram_inv(clk_mux_size3_32_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	clk_mux_size3 mux_bottom_track_67 (
		.in({chany_top_in[33], chanx_right_in[33], chanx_left_in[33]}),
		.sram(clk_mux_size3_33_sram[0:1]),
		.sram_inv(clk_mux_size3_33_sram_inv[0:1]),
		.out(chany_bottom_out[33]));

	clk_mux_size3 mux_bottom_track_69 (
		.in({chany_top_in[34], chanx_right_in[34], chanx_left_in[34]}),
		.sram(clk_mux_size3_34_sram[0:1]),
		.sram_inv(clk_mux_size3_34_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	clk_mux_size3 mux_bottom_track_71 (
		.in({chany_top_in[35], chanx_right_in[35], chanx_left_in[35]}),
		.sram(clk_mux_size3_35_sram[0:1]),
		.sram_inv(clk_mux_size3_35_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	clk_mux_size3 mux_bottom_track_73 (
		.in({chany_top_in[36], chanx_right_in[36], chanx_left_in[36]}),
		.sram(clk_mux_size3_36_sram[0:1]),
		.sram_inv(clk_mux_size3_36_sram_inv[0:1]),
		.out(chany_bottom_out[36]));

	clk_mux_size3 mux_bottom_track_75 (
		.in({chany_top_in[37], chanx_right_in[37], chanx_left_in[37]}),
		.sram(clk_mux_size3_37_sram[0:1]),
		.sram_inv(clk_mux_size3_37_sram_inv[0:1]),
		.out(chany_bottom_out[37]));

	clk_mux_size3 mux_bottom_track_77 (
		.in({chany_top_in[38], chanx_right_in[38], chanx_left_in[38]}),
		.sram(clk_mux_size3_38_sram[0:1]),
		.sram_inv(clk_mux_size3_38_sram_inv[0:1]),
		.out(chany_bottom_out[38]));

	clk_mux_size3 mux_bottom_track_79 (
		.in({chany_top_in[39], chanx_right_in[39], chanx_left_in[39]}),
		.sram(clk_mux_size3_39_sram[0:1]),
		.sram_inv(clk_mux_size3_39_sram_inv[0:1]),
		.out(chany_bottom_out[39]));

	clk_mux_size3 mux_bottom_track_81 (
		.in({chany_top_in[40], chanx_right_in[40], chanx_left_in[40]}),
		.sram(clk_mux_size3_40_sram[0:1]),
		.sram_inv(clk_mux_size3_40_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	clk_mux_size3 mux_bottom_track_83 (
		.in({chany_top_in[41], chanx_right_in[41], chanx_left_in[41]}),
		.sram(clk_mux_size3_41_sram[0:1]),
		.sram_inv(clk_mux_size3_41_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	clk_mux_size3 mux_bottom_track_85 (
		.in({chany_top_in[42], chanx_right_in[42], chanx_left_in[42]}),
		.sram(clk_mux_size3_42_sram[0:1]),
		.sram_inv(clk_mux_size3_42_sram_inv[0:1]),
		.out(chany_bottom_out[42]));

	clk_mux_size3 mux_bottom_track_87 (
		.in({chany_top_in[43], chanx_right_in[43], chanx_left_in[43]}),
		.sram(clk_mux_size3_43_sram[0:1]),
		.sram_inv(clk_mux_size3_43_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	clk_mux_size3 mux_bottom_track_89 (
		.in({chany_top_in[44], chanx_right_in[44], chanx_left_in[44]}),
		.sram(clk_mux_size3_44_sram[0:1]),
		.sram_inv(clk_mux_size3_44_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	clk_mux_size3 mux_bottom_track_91 (
		.in({chany_top_in[45], chanx_right_in[45], chanx_left_in[45]}),
		.sram(clk_mux_size3_45_sram[0:1]),
		.sram_inv(clk_mux_size3_45_sram_inv[0:1]),
		.out(chany_bottom_out[45]));

	clk_mux_size3 mux_bottom_track_93 (
		.in({chany_top_in[46], chanx_right_in[46], chanx_left_in[46]}),
		.sram(clk_mux_size3_46_sram[0:1]),
		.sram_inv(clk_mux_size3_46_sram_inv[0:1]),
		.out(chany_bottom_out[46]));

	clk_mux_size3 mux_bottom_track_95 (
		.in({chany_top_in[47], chanx_right_in[47], chanx_left_in[47]}),
		.sram(clk_mux_size3_47_sram[0:1]),
		.sram_inv(clk_mux_size3_47_sram_inv[0:1]),
		.out(chany_bottom_out[47]));

	clk_mux_size3 mux_bottom_track_97 (
		.in({chany_top_in[48], chanx_right_in[48], chanx_left_in[48]}),
		.sram(clk_mux_size3_48_sram[0:1]),
		.sram_inv(clk_mux_size3_48_sram_inv[0:1]),
		.out(chany_bottom_out[48]));

	clk_mux_size3 mux_bottom_track_99 (
		.in({chany_top_in[49], chanx_right_in[49], chanx_left_in[49]}),
		.sram(clk_mux_size3_49_sram[0:1]),
		.sram_inv(clk_mux_size3_49_sram_inv[0:1]),
		.out(chany_bottom_out[49]));

	clk_mux_size3 mux_bottom_track_101 (
		.in({chany_top_in[50], chanx_right_in[50], chanx_left_in[50]}),
		.sram(clk_mux_size3_50_sram[0:1]),
		.sram_inv(clk_mux_size3_50_sram_inv[0:1]),
		.out(chany_bottom_out[50]));

	clk_mux_size3 mux_bottom_track_103 (
		.in({chany_top_in[51], chanx_right_in[51], chanx_left_in[51]}),
		.sram(clk_mux_size3_51_sram[0:1]),
		.sram_inv(clk_mux_size3_51_sram_inv[0:1]),
		.out(chany_bottom_out[51]));

	clk_mux_size3 mux_bottom_track_105 (
		.in({chany_top_in[52], chanx_right_in[52], chanx_left_in[52]}),
		.sram(clk_mux_size3_52_sram[0:1]),
		.sram_inv(clk_mux_size3_52_sram_inv[0:1]),
		.out(chany_bottom_out[52]));

	clk_mux_size3 mux_bottom_track_107 (
		.in({chany_top_in[53], chanx_right_in[53], chanx_left_in[53]}),
		.sram(clk_mux_size3_53_sram[0:1]),
		.sram_inv(clk_mux_size3_53_sram_inv[0:1]),
		.out(chany_bottom_out[53]));

	clk_mux_size3 mux_bottom_track_109 (
		.in({chany_top_in[54], chanx_right_in[54], chanx_left_in[54]}),
		.sram(clk_mux_size3_54_sram[0:1]),
		.sram_inv(clk_mux_size3_54_sram_inv[0:1]),
		.out(chany_bottom_out[54]));

	clk_mux_size3 mux_bottom_track_111 (
		.in({chany_top_in[55], chanx_right_in[55], chanx_left_in[55]}),
		.sram(clk_mux_size3_55_sram[0:1]),
		.sram_inv(clk_mux_size3_55_sram_inv[0:1]),
		.out(chany_bottom_out[55]));

	clk_mux_size3 mux_bottom_track_113 (
		.in({chany_top_in[56], chanx_right_in[56], chanx_left_in[56]}),
		.sram(clk_mux_size3_56_sram[0:1]),
		.sram_inv(clk_mux_size3_56_sram_inv[0:1]),
		.out(chany_bottom_out[56]));

	clk_mux_size3 mux_bottom_track_115 (
		.in({chany_top_in[57], chanx_right_in[57], chanx_left_in[57]}),
		.sram(clk_mux_size3_57_sram[0:1]),
		.sram_inv(clk_mux_size3_57_sram_inv[0:1]),
		.out(chany_bottom_out[57]));

	clk_mux_size3 mux_bottom_track_117 (
		.in({chany_top_in[58], chanx_right_in[58], chanx_left_in[58]}),
		.sram(clk_mux_size3_58_sram[0:1]),
		.sram_inv(clk_mux_size3_58_sram_inv[0:1]),
		.out(chany_bottom_out[58]));

	clk_mux_size3 mux_bottom_track_119 (
		.in({chany_top_in[59], chanx_right_in[59], chanx_left_in[59]}),
		.sram(clk_mux_size3_59_sram[0:1]),
		.sram_inv(clk_mux_size3_59_sram_inv[0:1]),
		.out(chany_bottom_out[59]));

	clk_mux_size3 mux_bottom_track_121 (
		.in({chany_top_in[60], chanx_right_in[60], chanx_left_in[60]}),
		.sram(clk_mux_size3_60_sram[0:1]),
		.sram_inv(clk_mux_size3_60_sram_inv[0:1]),
		.out(chany_bottom_out[60]));

	clk_mux_size3 mux_bottom_track_123 (
		.in({chany_top_in[61], chanx_right_in[61], chanx_left_in[61]}),
		.sram(clk_mux_size3_61_sram[0:1]),
		.sram_inv(clk_mux_size3_61_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	clk_mux_size3 mux_bottom_track_125 (
		.in({chany_top_in[62], chanx_right_in[62], chanx_left_in[62]}),
		.sram(clk_mux_size3_62_sram[0:1]),
		.sram_inv(clk_mux_size3_62_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	clk_mux_size3 mux_bottom_track_127 (
		.in({chany_top_in[63], chanx_right_in[63], chanx_left_in[63]}),
		.sram(clk_mux_size3_63_sram[0:1]),
		.sram_inv(clk_mux_size3_63_sram_inv[0:1]),
		.out(chany_bottom_out[63]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_64 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[54:55]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[54:55]),
		.mem_out(clk_mux_size3_0_sram[0:1]),
		.mem_outb(clk_mux_size3_0_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_66 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[56:57]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[56:57]),
		.mem_out(clk_mux_size3_1_sram[0:1]),
		.mem_outb(clk_mux_size3_1_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_68 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[58:59]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[58:59]),
		.mem_out(clk_mux_size3_2_sram[0:1]),
		.mem_outb(clk_mux_size3_2_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_70 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[60:61]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[60:61]),
		.mem_out(clk_mux_size3_3_sram[0:1]),
		.mem_outb(clk_mux_size3_3_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_72 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[62:63]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[62:63]),
		.mem_out(clk_mux_size3_4_sram[0:1]),
		.mem_outb(clk_mux_size3_4_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_74 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[64:65]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[64:65]),
		.mem_out(clk_mux_size3_5_sram[0:1]),
		.mem_outb(clk_mux_size3_5_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_76 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[66:67]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[66:67]),
		.mem_out(clk_mux_size3_6_sram[0:1]),
		.mem_outb(clk_mux_size3_6_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_78 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[68:69]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[68:69]),
		.mem_out(clk_mux_size3_7_sram[0:1]),
		.mem_outb(clk_mux_size3_7_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_80 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[70:71]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[70:71]),
		.mem_out(clk_mux_size3_8_sram[0:1]),
		.mem_outb(clk_mux_size3_8_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_82 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[72:73]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[72:73]),
		.mem_out(clk_mux_size3_9_sram[0:1]),
		.mem_outb(clk_mux_size3_9_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_84 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[74:75]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[74:75]),
		.mem_out(clk_mux_size3_10_sram[0:1]),
		.mem_outb(clk_mux_size3_10_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_86 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[76:77]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[76:77]),
		.mem_out(clk_mux_size3_11_sram[0:1]),
		.mem_outb(clk_mux_size3_11_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_88 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[78:79]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[78:79]),
		.mem_out(clk_mux_size3_12_sram[0:1]),
		.mem_outb(clk_mux_size3_12_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_90 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[80:81]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[80:81]),
		.mem_out(clk_mux_size3_13_sram[0:1]),
		.mem_outb(clk_mux_size3_13_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_92 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[82:83]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[82:83]),
		.mem_out(clk_mux_size3_14_sram[0:1]),
		.mem_outb(clk_mux_size3_14_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_94 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[84:85]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[84:85]),
		.mem_out(clk_mux_size3_15_sram[0:1]),
		.mem_outb(clk_mux_size3_15_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_96 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[86:87]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[86:87]),
		.mem_out(clk_mux_size3_16_sram[0:1]),
		.mem_outb(clk_mux_size3_16_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_98 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[88:89]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[88:89]),
		.mem_out(clk_mux_size3_17_sram[0:1]),
		.mem_outb(clk_mux_size3_17_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_100 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[90:91]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[90:91]),
		.mem_out(clk_mux_size3_18_sram[0:1]),
		.mem_outb(clk_mux_size3_18_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_102 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[92:93]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[92:93]),
		.mem_out(clk_mux_size3_19_sram[0:1]),
		.mem_outb(clk_mux_size3_19_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_104 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[94:95]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[94:95]),
		.mem_out(clk_mux_size3_20_sram[0:1]),
		.mem_outb(clk_mux_size3_20_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_106 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[96:97]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[96:97]),
		.mem_out(clk_mux_size3_21_sram[0:1]),
		.mem_outb(clk_mux_size3_21_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_108 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[98:99]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[98:99]),
		.mem_out(clk_mux_size3_22_sram[0:1]),
		.mem_outb(clk_mux_size3_22_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_110 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[100:101]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[100:101]),
		.mem_out(clk_mux_size3_23_sram[0:1]),
		.mem_outb(clk_mux_size3_23_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_112 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[102:103]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[102:103]),
		.mem_out(clk_mux_size3_24_sram[0:1]),
		.mem_outb(clk_mux_size3_24_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_114 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[104:105]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[104:105]),
		.mem_out(clk_mux_size3_25_sram[0:1]),
		.mem_outb(clk_mux_size3_25_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_116 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[106:107]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[106:107]),
		.mem_out(clk_mux_size3_26_sram[0:1]),
		.mem_outb(clk_mux_size3_26_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_118 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[108:109]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[108:109]),
		.mem_out(clk_mux_size3_27_sram[0:1]),
		.mem_outb(clk_mux_size3_27_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_120 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[110:111]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[110:111]),
		.mem_out(clk_mux_size3_28_sram[0:1]),
		.mem_outb(clk_mux_size3_28_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_122 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[112:113]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[112:113]),
		.mem_out(clk_mux_size3_29_sram[0:1]),
		.mem_outb(clk_mux_size3_29_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_124 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[114:115]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[114:115]),
		.mem_out(clk_mux_size3_30_sram[0:1]),
		.mem_outb(clk_mux_size3_30_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_126 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[116:117]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[116:117]),
		.mem_out(clk_mux_size3_31_sram[0:1]),
		.mem_outb(clk_mux_size3_31_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_65 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[224:225]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[224:225]),
		.mem_out(clk_mux_size3_32_sram[0:1]),
		.mem_outb(clk_mux_size3_32_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_67 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[226:227]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[226:227]),
		.mem_out(clk_mux_size3_33_sram[0:1]),
		.mem_outb(clk_mux_size3_33_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_69 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[228:229]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[228:229]),
		.mem_out(clk_mux_size3_34_sram[0:1]),
		.mem_outb(clk_mux_size3_34_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_71 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[230:231]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[230:231]),
		.mem_out(clk_mux_size3_35_sram[0:1]),
		.mem_outb(clk_mux_size3_35_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_73 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[232:233]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[232:233]),
		.mem_out(clk_mux_size3_36_sram[0:1]),
		.mem_outb(clk_mux_size3_36_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_75 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[234:235]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[234:235]),
		.mem_out(clk_mux_size3_37_sram[0:1]),
		.mem_outb(clk_mux_size3_37_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_77 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[236:237]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[236:237]),
		.mem_out(clk_mux_size3_38_sram[0:1]),
		.mem_outb(clk_mux_size3_38_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_79 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[238:239]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[238:239]),
		.mem_out(clk_mux_size3_39_sram[0:1]),
		.mem_outb(clk_mux_size3_39_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_81 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[240:241]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[240:241]),
		.mem_out(clk_mux_size3_40_sram[0:1]),
		.mem_outb(clk_mux_size3_40_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_83 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[242:243]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[242:243]),
		.mem_out(clk_mux_size3_41_sram[0:1]),
		.mem_outb(clk_mux_size3_41_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_85 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[244:245]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[244:245]),
		.mem_out(clk_mux_size3_42_sram[0:1]),
		.mem_outb(clk_mux_size3_42_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_87 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[246:247]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[246:247]),
		.mem_out(clk_mux_size3_43_sram[0:1]),
		.mem_outb(clk_mux_size3_43_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_89 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[248:249]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[248:249]),
		.mem_out(clk_mux_size3_44_sram[0:1]),
		.mem_outb(clk_mux_size3_44_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_91 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[250:251]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[250:251]),
		.mem_out(clk_mux_size3_45_sram[0:1]),
		.mem_outb(clk_mux_size3_45_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_93 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[252:253]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[252:253]),
		.mem_out(clk_mux_size3_46_sram[0:1]),
		.mem_outb(clk_mux_size3_46_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_95 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[254:255]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[254:255]),
		.mem_out(clk_mux_size3_47_sram[0:1]),
		.mem_outb(clk_mux_size3_47_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_97 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[256:257]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[256:257]),
		.mem_out(clk_mux_size3_48_sram[0:1]),
		.mem_outb(clk_mux_size3_48_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_99 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[258:259]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[258:259]),
		.mem_out(clk_mux_size3_49_sram[0:1]),
		.mem_outb(clk_mux_size3_49_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_101 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[260:261]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[260:261]),
		.mem_out(clk_mux_size3_50_sram[0:1]),
		.mem_outb(clk_mux_size3_50_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_103 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[262:263]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[262:263]),
		.mem_out(clk_mux_size3_51_sram[0:1]),
		.mem_outb(clk_mux_size3_51_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_105 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[264:265]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[264:265]),
		.mem_out(clk_mux_size3_52_sram[0:1]),
		.mem_outb(clk_mux_size3_52_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_107 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[266:267]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[266:267]),
		.mem_out(clk_mux_size3_53_sram[0:1]),
		.mem_outb(clk_mux_size3_53_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_109 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[268:269]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[268:269]),
		.mem_out(clk_mux_size3_54_sram[0:1]),
		.mem_outb(clk_mux_size3_54_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_111 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[270:271]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[270:271]),
		.mem_out(clk_mux_size3_55_sram[0:1]),
		.mem_outb(clk_mux_size3_55_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_113 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[272:273]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[272:273]),
		.mem_out(clk_mux_size3_56_sram[0:1]),
		.mem_outb(clk_mux_size3_56_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_115 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[274:275]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[274:275]),
		.mem_out(clk_mux_size3_57_sram[0:1]),
		.mem_outb(clk_mux_size3_57_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_117 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[276:277]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[276:277]),
		.mem_out(clk_mux_size3_58_sram[0:1]),
		.mem_outb(clk_mux_size3_58_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_119 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[278:279]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[278:279]),
		.mem_out(clk_mux_size3_59_sram[0:1]),
		.mem_outb(clk_mux_size3_59_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_121 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[280:281]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[280:281]),
		.mem_out(clk_mux_size3_60_sram[0:1]),
		.mem_outb(clk_mux_size3_60_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_123 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[282:283]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[282:283]),
		.mem_out(clk_mux_size3_61_sram[0:1]),
		.mem_outb(clk_mux_size3_61_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_125 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[284:285]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[284:285]),
		.mem_out(clk_mux_size3_62_sram[0:1]),
		.mem_outb(clk_mux_size3_62_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_127 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[286:287]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[286:287]),
		.mem_out(clk_mux_size3_63_sram[0:1]),
		.mem_outb(clk_mux_size3_63_sram_inv[0:1]));

	sb_mux_size11 mux_right_track_0 (
		.in({chany_top_in[6], chany_top_in[26], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[6], chany_bottom_in[26:27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[0]}),
		.sram(sb_mux_size11_0_sram[0:3]),
		.sram_inv(sb_mux_size11_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	sb_mux_size11 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[8], chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[8], chany_bottom_in[23], chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[1]}),
		.sram(sb_mux_size11_1_sram[0:3]),
		.sram_inv(sb_mux_size11_1_sram_inv[0:3]),
		.out(chanx_right_out[1]));

	sb_mux_size11 mux_right_track_12 (
		.in({chany_top_in[5], chany_top_in[16], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chany_bottom_in[7], chany_bottom_in[16], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[7]}),
		.sram(sb_mux_size11_2_sram[0:3]),
		.sram_inv(sb_mux_size11_2_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	sb_mux_size11 mux_right_track_16 (
		.in({chany_top_in[7], chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chany_bottom_in[5], chany_bottom_in[17], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[9]}),
		.sram(sb_mux_size11_3_sram[0:3]),
		.sram_inv(sb_mux_size11_3_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	sb_mux_size11 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[6], chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[0], chany_bottom_in[6], chany_bottom_in[26], chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_}),
		.sram(sb_mux_size11_4_sram[0:3]),
		.sram_inv(sb_mux_size11_4_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	sb_mux_size11 mux_left_track_3 (
		.in({chany_top_in[8], chany_top_in[28], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[1], chany_bottom_in[0], chany_bottom_in[8], chany_bottom_in[28], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_}),
		.sram(sb_mux_size11_5_sram[0:3]),
		.sram_inv(sb_mux_size11_5_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	sb_mux_size11 mux_left_track_13 (
		.in({chany_top_in[11], chany_top_in[16], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[7], chany_bottom_in[5], chany_bottom_in[16], left_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_}),
		.sram(sb_mux_size11_6_sram[0:3]),
		.sram_inv(sb_mux_size11_6_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	sb_mux_size11 mux_left_track_17 (
		.in({chany_top_in[9], chany_top_in[17], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[9], chany_bottom_in[7], chany_bottom_in[17], left_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_}),
		.sram(sb_mux_size11_7_sram[0:3]),
		.sram_inv(sb_mux_size11_7_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_right_track_0 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[118:121]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[118:121]),
		.mem_out(sb_mux_size11_0_sram[0:3]),
		.mem_outb(sb_mux_size11_0_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_right_track_2 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[122:125]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[122:125]),
		.mem_out(sb_mux_size11_1_sram[0:3]),
		.mem_outb(sb_mux_size11_1_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_right_track_12 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[140:143]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[140:143]),
		.mem_out(sb_mux_size11_2_sram[0:3]),
		.mem_outb(sb_mux_size11_2_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_right_track_16 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[144:147]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[144:147]),
		.mem_out(sb_mux_size11_3_sram[0:3]),
		.mem_outb(sb_mux_size11_3_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_left_track_1 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[288:291]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[288:291]),
		.mem_out(sb_mux_size11_4_sram[0:3]),
		.mem_outb(sb_mux_size11_4_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_left_track_3 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[292:295]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[292:295]),
		.mem_out(sb_mux_size11_5_sram[0:3]),
		.mem_outb(sb_mux_size11_5_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_left_track_13 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[310:313]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[310:313]),
		.mem_out(sb_mux_size11_6_sram[0:3]),
		.mem_outb(sb_mux_size11_6_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_left_track_17 (
		.feedthrough_mem_in(sb_6__config_group_mem_size340_0_mem_out[314:317]),
		.feedthrough_mem_inb(sb_6__config_group_mem_size340_0_mem_outb[314:317]),
		.mem_out(sb_mux_size11_7_sram[0:3]),
		.mem_outb(sb_mux_size11_7_sram_inv[0:3]));

	sb_6__config_group_mem_size340 sb_6__config_group_mem_size340 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.mem_out(sb_6__config_group_mem_size340_0_mem_out[0:339]),
		.mem_outb(sb_6__config_group_mem_size340_0_mem_outb[0:339]),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for sb_6_ -----



