//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Connection Blocks[0][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for cby_1_ -----
module cby_1_(config_enable,
              prog_reset,
              prog_clk,
              chany_bottom_in,
              chany_top_in,
              ccff_head,
              chany_bottom_out,
              chany_top_out,
              left_grid_right_width_0_height_0_subtile_0__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_0__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_1__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_1__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_2__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_2__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_3__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_3__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_4__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_4__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_5__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_5__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_6__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_6__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_7__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_7__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_8__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_8__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_9__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_9__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_10__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_10__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_11__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_11__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_12__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_12__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_13__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_13__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_14__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_14__pin_clk_0_,
              left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_,
              left_grid_right_width_0_height_0_subtile_15__pin_reset_0_,
              left_grid_right_width_0_height_0_subtile_15__pin_clk_0_,
              ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:63] chany_bottom_in;
//----- INPUT PORTS -----
input [0:63] chany_top_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:63] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:63] chany_top_out;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_1__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_1__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_2__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_2__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_3__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_3__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_4__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_4__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_5__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_5__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_6__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_6__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_7__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_7__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_8__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_8__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_9__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_9__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_10__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_10__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_11__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_11__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_12__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_12__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_13__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_13__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_14__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_14__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_15__pin_reset_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_15__pin_clk_0_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:4] cb_mux_size16_0_sram;
wire [0:4] cb_mux_size16_0_sram_inv;
wire [0:4] cb_mux_size16_10_sram;
wire [0:4] cb_mux_size16_10_sram_inv;
wire [0:4] cb_mux_size16_11_sram;
wire [0:4] cb_mux_size16_11_sram_inv;
wire [0:4] cb_mux_size16_12_sram;
wire [0:4] cb_mux_size16_12_sram_inv;
wire [0:4] cb_mux_size16_13_sram;
wire [0:4] cb_mux_size16_13_sram_inv;
wire [0:4] cb_mux_size16_14_sram;
wire [0:4] cb_mux_size16_14_sram_inv;
wire [0:4] cb_mux_size16_15_sram;
wire [0:4] cb_mux_size16_15_sram_inv;
wire [0:4] cb_mux_size16_1_sram;
wire [0:4] cb_mux_size16_1_sram_inv;
wire [0:4] cb_mux_size16_2_sram;
wire [0:4] cb_mux_size16_2_sram_inv;
wire [0:4] cb_mux_size16_3_sram;
wire [0:4] cb_mux_size16_3_sram_inv;
wire [0:4] cb_mux_size16_4_sram;
wire [0:4] cb_mux_size16_4_sram_inv;
wire [0:4] cb_mux_size16_5_sram;
wire [0:4] cb_mux_size16_5_sram_inv;
wire [0:4] cb_mux_size16_6_sram;
wire [0:4] cb_mux_size16_6_sram_inv;
wire [0:4] cb_mux_size16_7_sram;
wire [0:4] cb_mux_size16_7_sram_inv;
wire [0:4] cb_mux_size16_8_sram;
wire [0:4] cb_mux_size16_8_sram_inv;
wire [0:4] cb_mux_size16_9_sram;
wire [0:4] cb_mux_size16_9_sram_inv;
wire [0:5] cb_mux_size48_0_sram;
wire [0:5] cb_mux_size48_0_sram_inv;
wire [0:5] cb_mux_size48_10_sram;
wire [0:5] cb_mux_size48_10_sram_inv;
wire [0:5] cb_mux_size48_11_sram;
wire [0:5] cb_mux_size48_11_sram_inv;
wire [0:5] cb_mux_size48_12_sram;
wire [0:5] cb_mux_size48_12_sram_inv;
wire [0:5] cb_mux_size48_13_sram;
wire [0:5] cb_mux_size48_13_sram_inv;
wire [0:5] cb_mux_size48_14_sram;
wire [0:5] cb_mux_size48_14_sram_inv;
wire [0:5] cb_mux_size48_15_sram;
wire [0:5] cb_mux_size48_15_sram_inv;
wire [0:5] cb_mux_size48_1_sram;
wire [0:5] cb_mux_size48_1_sram_inv;
wire [0:5] cb_mux_size48_2_sram;
wire [0:5] cb_mux_size48_2_sram_inv;
wire [0:5] cb_mux_size48_3_sram;
wire [0:5] cb_mux_size48_3_sram_inv;
wire [0:5] cb_mux_size48_4_sram;
wire [0:5] cb_mux_size48_4_sram_inv;
wire [0:5] cb_mux_size48_5_sram;
wire [0:5] cb_mux_size48_5_sram_inv;
wire [0:5] cb_mux_size48_6_sram;
wire [0:5] cb_mux_size48_6_sram_inv;
wire [0:5] cb_mux_size48_7_sram;
wire [0:5] cb_mux_size48_7_sram_inv;
wire [0:5] cb_mux_size48_8_sram;
wire [0:5] cb_mux_size48_8_sram_inv;
wire [0:5] cb_mux_size48_9_sram;
wire [0:5] cb_mux_size48_9_sram_inv;
wire [0:5] cb_mux_size56_0_sram;
wire [0:5] cb_mux_size56_0_sram_inv;
wire [0:5] cb_mux_size56_1_sram;
wire [0:5] cb_mux_size56_1_sram_inv;
wire [0:5] cb_mux_size56_2_sram;
wire [0:5] cb_mux_size56_2_sram_inv;
wire [0:5] cb_mux_size56_3_sram;
wire [0:5] cb_mux_size56_3_sram_inv;
wire [0:5] cb_mux_size56_4_sram;
wire [0:5] cb_mux_size56_4_sram_inv;
wire [0:5] cb_mux_size56_5_sram;
wire [0:5] cb_mux_size56_5_sram_inv;
wire [0:5] cb_mux_size56_6_sram;
wire [0:5] cb_mux_size56_6_sram_inv;
wire [0:5] cb_mux_size56_7_sram;
wire [0:5] cb_mux_size56_7_sram_inv;
wire [0:223] cby_1__config_group_mem_size224_0_mem_out;
wire [0:223] cby_1__config_group_mem_size224_0_mem_outb;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[0] = chany_bottom_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[4] = chany_bottom_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chany_bottom_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[12] = chany_bottom_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[16] = chany_bottom_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[20] = chany_bottom_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[24] = chany_bottom_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[28] = chany_bottom_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[32] = chany_bottom_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[36] = chany_bottom_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[40] = chany_bottom_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chany_bottom_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[48] = chany_bottom_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[52] = chany_bottom_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[56] = chany_bottom_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chany_bottom_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[0] = chany_top_in[0];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[1];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[2];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[3];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[4] = chany_top_in[4];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[5];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[6];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[7];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[8] = chany_top_in[8];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[9];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[10];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[11];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[12] = chany_top_in[12];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[13];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[14];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[15];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[16] = chany_top_in[16];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[17];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[18];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[19];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[20] = chany_top_in[20];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[21];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[22];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[23];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[24] = chany_top_in[24];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[25];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[26];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[27];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[28] = chany_top_in[28];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[29];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[30];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[31];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[32] = chany_top_in[32];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[33];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[34];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[35];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[36] = chany_top_in[36];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[37];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[38];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[39];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[40] = chany_top_in[40];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[41];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[42];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[43];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[44] = chany_top_in[44];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[45];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[46];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[47];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[48] = chany_top_in[48];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[49];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[50];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[51];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[52] = chany_top_in[52];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[53];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[54];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[55];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[56] = chany_top_in[56];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[57];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[58];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[59];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[60] = chany_top_in[60];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[61];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[62];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[63];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size48 mux_right_ipin_0 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_0_sram[0:5]),
		.sram_inv(cb_mux_size48_0_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_2 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_1_sram[0:5]),
		.sram_inv(cb_mux_size48_1_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_1__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_4 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_2_sram[0:5]),
		.sram_inv(cb_mux_size48_2_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_2__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_6 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_3_sram[0:5]),
		.sram_inv(cb_mux_size48_3_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_3__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_8 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_4_sram[0:5]),
		.sram_inv(cb_mux_size48_4_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_4__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_10 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_5_sram[0:5]),
		.sram_inv(cb_mux_size48_5_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_5__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_12 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_6_sram[0:5]),
		.sram_inv(cb_mux_size48_6_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_6__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_14 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_7_sram[0:5]),
		.sram_inv(cb_mux_size48_7_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_7__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_17 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_8_sram[0:5]),
		.sram_inv(cb_mux_size48_8_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_8__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_20 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_9_sram[0:5]),
		.sram_inv(cb_mux_size48_9_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_9__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_23 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_10_sram[0:5]),
		.sram_inv(cb_mux_size48_10_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_10__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_26 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_11_sram[0:5]),
		.sram_inv(cb_mux_size48_11_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_11__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_29 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_12_sram[0:5]),
		.sram_inv(cb_mux_size48_12_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_12__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_32 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_13_sram[0:5]),
		.sram_inv(cb_mux_size48_13_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_13__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_35 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_14_sram[0:5]),
		.sram_inv(cb_mux_size48_14_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_14__pin_reset_0_));

	cb_mux_size48 mux_right_ipin_38 (
		.in({chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size48_15_sram[0:5]),
		.sram_inv(cb_mux_size48_15_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_15__pin_reset_0_));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_0 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[0:5]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[0:5]),
		.mem_out(cb_mux_size48_0_sram[0:5]),
		.mem_outb(cb_mux_size48_0_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_2 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[11:16]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[11:16]),
		.mem_out(cb_mux_size48_1_sram[0:5]),
		.mem_outb(cb_mux_size48_1_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_4 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[22:27]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[22:27]),
		.mem_out(cb_mux_size48_2_sram[0:5]),
		.mem_outb(cb_mux_size48_2_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_6 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[33:38]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[33:38]),
		.mem_out(cb_mux_size48_3_sram[0:5]),
		.mem_outb(cb_mux_size48_3_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_8 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[44:49]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[44:49]),
		.mem_out(cb_mux_size48_4_sram[0:5]),
		.mem_outb(cb_mux_size48_4_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_10 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[55:60]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[55:60]),
		.mem_out(cb_mux_size48_5_sram[0:5]),
		.mem_outb(cb_mux_size48_5_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_12 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[66:71]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[66:71]),
		.mem_out(cb_mux_size48_6_sram[0:5]),
		.mem_outb(cb_mux_size48_6_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_14 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[77:82]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[77:82]),
		.mem_out(cb_mux_size48_7_sram[0:5]),
		.mem_outb(cb_mux_size48_7_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_17 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[94:99]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[94:99]),
		.mem_out(cb_mux_size48_8_sram[0:5]),
		.mem_outb(cb_mux_size48_8_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_20 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[111:116]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[111:116]),
		.mem_out(cb_mux_size48_9_sram[0:5]),
		.mem_outb(cb_mux_size48_9_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_23 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[128:133]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[128:133]),
		.mem_out(cb_mux_size48_10_sram[0:5]),
		.mem_outb(cb_mux_size48_10_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_26 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[145:150]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[145:150]),
		.mem_out(cb_mux_size48_11_sram[0:5]),
		.mem_outb(cb_mux_size48_11_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_29 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[162:167]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[162:167]),
		.mem_out(cb_mux_size48_12_sram[0:5]),
		.mem_outb(cb_mux_size48_12_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_32 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[179:184]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[179:184]),
		.mem_out(cb_mux_size48_13_sram[0:5]),
		.mem_outb(cb_mux_size48_13_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_35 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[196:201]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[196:201]),
		.mem_out(cb_mux_size48_14_sram[0:5]),
		.mem_outb(cb_mux_size48_14_sram_inv[0:5]));

	cb_mux_size48_feedthrough_mem feedthrough_mem_right_ipin_38 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[213:218]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[213:218]),
		.mem_out(cb_mux_size48_15_sram[0:5]),
		.mem_outb(cb_mux_size48_15_sram_inv[0:5]));

	cb_mux_size16 mux_right_ipin_1 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_0_sram[0:4]),
		.sram_inv(cb_mux_size16_0_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_3 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_1_sram[0:4]),
		.sram_inv(cb_mux_size16_1_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_1__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_5 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_2_sram[0:4]),
		.sram_inv(cb_mux_size16_2_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_2__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_7 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_3_sram[0:4]),
		.sram_inv(cb_mux_size16_3_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_3__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_9 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_4_sram[0:4]),
		.sram_inv(cb_mux_size16_4_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_4__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_11 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_5_sram[0:4]),
		.sram_inv(cb_mux_size16_5_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_5__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_13 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_6_sram[0:4]),
		.sram_inv(cb_mux_size16_6_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_6__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_15 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_7_sram[0:4]),
		.sram_inv(cb_mux_size16_7_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_7__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_18 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_8_sram[0:4]),
		.sram_inv(cb_mux_size16_8_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_8__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_21 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_9_sram[0:4]),
		.sram_inv(cb_mux_size16_9_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_9__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_24 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_10_sram[0:4]),
		.sram_inv(cb_mux_size16_10_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_10__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_27 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_11_sram[0:4]),
		.sram_inv(cb_mux_size16_11_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_11__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_30 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_12_sram[0:4]),
		.sram_inv(cb_mux_size16_12_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_12__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_33 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_13_sram[0:4]),
		.sram_inv(cb_mux_size16_13_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_13__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_36 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_14_sram[0:4]),
		.sram_inv(cb_mux_size16_14_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_14__pin_clk_0_));

	cb_mux_size16 mux_right_ipin_39 (
		.in({chany_bottom_in[32], chany_top_in[32], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[39], chany_top_in[39]}),
		.sram(cb_mux_size16_15_sram[0:4]),
		.sram_inv(cb_mux_size16_15_sram_inv[0:4]),
		.out(left_grid_right_width_0_height_0_subtile_15__pin_clk_0_));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_1 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[6:10]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[6:10]),
		.mem_out(cb_mux_size16_0_sram[0:4]),
		.mem_outb(cb_mux_size16_0_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_3 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[17:21]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[17:21]),
		.mem_out(cb_mux_size16_1_sram[0:4]),
		.mem_outb(cb_mux_size16_1_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_5 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[28:32]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[28:32]),
		.mem_out(cb_mux_size16_2_sram[0:4]),
		.mem_outb(cb_mux_size16_2_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_7 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[39:43]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[39:43]),
		.mem_out(cb_mux_size16_3_sram[0:4]),
		.mem_outb(cb_mux_size16_3_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_9 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[50:54]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[50:54]),
		.mem_out(cb_mux_size16_4_sram[0:4]),
		.mem_outb(cb_mux_size16_4_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_11 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[61:65]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[61:65]),
		.mem_out(cb_mux_size16_5_sram[0:4]),
		.mem_outb(cb_mux_size16_5_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_13 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[72:76]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[72:76]),
		.mem_out(cb_mux_size16_6_sram[0:4]),
		.mem_outb(cb_mux_size16_6_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_15 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[83:87]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[83:87]),
		.mem_out(cb_mux_size16_7_sram[0:4]),
		.mem_outb(cb_mux_size16_7_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_18 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[100:104]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[100:104]),
		.mem_out(cb_mux_size16_8_sram[0:4]),
		.mem_outb(cb_mux_size16_8_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_21 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[117:121]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[117:121]),
		.mem_out(cb_mux_size16_9_sram[0:4]),
		.mem_outb(cb_mux_size16_9_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_24 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[134:138]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[134:138]),
		.mem_out(cb_mux_size16_10_sram[0:4]),
		.mem_outb(cb_mux_size16_10_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_27 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[151:155]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[151:155]),
		.mem_out(cb_mux_size16_11_sram[0:4]),
		.mem_outb(cb_mux_size16_11_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_30 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[168:172]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[168:172]),
		.mem_out(cb_mux_size16_12_sram[0:4]),
		.mem_outb(cb_mux_size16_12_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_33 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[185:189]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[185:189]),
		.mem_out(cb_mux_size16_13_sram[0:4]),
		.mem_outb(cb_mux_size16_13_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_36 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[202:206]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[202:206]),
		.mem_out(cb_mux_size16_14_sram[0:4]),
		.mem_outb(cb_mux_size16_14_sram_inv[0:4]));

	cb_mux_size16_feedthrough_mem feedthrough_mem_right_ipin_39 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[219:223]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[219:223]),
		.mem_out(cb_mux_size16_15_sram[0:4]),
		.mem_outb(cb_mux_size16_15_sram_inv[0:4]));

	cb_mux_size56 mux_right_ipin_16 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_0_sram[0:5]),
		.sram_inv(cb_mux_size56_0_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_8__pin_f2a_i_0_));

	cb_mux_size56 mux_right_ipin_19 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_1_sram[0:5]),
		.sram_inv(cb_mux_size56_1_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_9__pin_f2a_i_0_));

	cb_mux_size56 mux_right_ipin_22 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_2_sram[0:5]),
		.sram_inv(cb_mux_size56_2_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_10__pin_f2a_i_0_));

	cb_mux_size56 mux_right_ipin_25 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_3_sram[0:5]),
		.sram_inv(cb_mux_size56_3_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_11__pin_f2a_i_0_));

	cb_mux_size56 mux_right_ipin_28 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_4_sram[0:5]),
		.sram_inv(cb_mux_size56_4_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_12__pin_f2a_i_0_));

	cb_mux_size56 mux_right_ipin_31 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_5_sram[0:5]),
		.sram_inv(cb_mux_size56_5_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_13__pin_f2a_i_0_));

	cb_mux_size56 mux_right_ipin_34 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_6_sram[0:5]),
		.sram_inv(cb_mux_size56_6_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_14__pin_f2a_i_0_));

	cb_mux_size56 mux_right_ipin_37 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[63], chany_top_in[63]}),
		.sram(cb_mux_size56_7_sram[0:5]),
		.sram_inv(cb_mux_size56_7_sram_inv[0:5]),
		.out(left_grid_right_width_0_height_0_subtile_15__pin_f2a_i_0_));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_16 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[88:93]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[88:93]),
		.mem_out(cb_mux_size56_0_sram[0:5]),
		.mem_outb(cb_mux_size56_0_sram_inv[0:5]));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_19 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[105:110]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[105:110]),
		.mem_out(cb_mux_size56_1_sram[0:5]),
		.mem_outb(cb_mux_size56_1_sram_inv[0:5]));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_22 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[122:127]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[122:127]),
		.mem_out(cb_mux_size56_2_sram[0:5]),
		.mem_outb(cb_mux_size56_2_sram_inv[0:5]));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_25 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[139:144]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[139:144]),
		.mem_out(cb_mux_size56_3_sram[0:5]),
		.mem_outb(cb_mux_size56_3_sram_inv[0:5]));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_28 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[156:161]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[156:161]),
		.mem_out(cb_mux_size56_4_sram[0:5]),
		.mem_outb(cb_mux_size56_4_sram_inv[0:5]));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_31 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[173:178]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[173:178]),
		.mem_out(cb_mux_size56_5_sram[0:5]),
		.mem_outb(cb_mux_size56_5_sram_inv[0:5]));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_34 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[190:195]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[190:195]),
		.mem_out(cb_mux_size56_6_sram[0:5]),
		.mem_outb(cb_mux_size56_6_sram_inv[0:5]));

	cb_mux_size56_feedthrough_mem feedthrough_mem_right_ipin_37 (
		.feedthrough_mem_in(cby_1__config_group_mem_size224_0_mem_out[207:212]),
		.feedthrough_mem_inb(cby_1__config_group_mem_size224_0_mem_outb[207:212]),
		.mem_out(cb_mux_size56_7_sram[0:5]),
		.mem_outb(cb_mux_size56_7_sram_inv[0:5]));

	cby_1__config_group_mem_size224 cby_1__config_group_mem_size224 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.mem_out(cby_1__config_group_mem_size224_0_mem_out[0:223]),
		.mem_outb(cby_1__config_group_mem_size224_0_mem_outb[0:223]),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for cby_1_ -----




