//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Wrapper Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for fpga_core -----
module fpga_core(clk,
                 reset,
                 prog_clk,
                 SE0,
                 SE1,
                 SC0,
                 SC1,
                 SR,
                 SE2,
                 config_enable,
                 prog_reset,
                 gfpga_pad_pinput_extmode_A2F,
                 gfpga_pad_pinput_dchain_extmode_A2F,
                 gfpga_pad_pinput_extmode_mode_o,
                 gfpga_pad_poutput_F2A,
                 gfpga_pad_mmffosc2cko_wrapper_C_O,
                 gfpga_pad_pinput_dchain_extmode_mode_o,
                 ccff_head,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:7] clk;
//----- GLOBAL PORTS -----
input [0:23] reset;
//----- GLOBAL PORTS -----
input [0:7] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] SE0;
//----- GLOBAL PORTS -----
input [0:0] SE1;
//----- GLOBAL PORTS -----
input [0:0] SC0;
//----- GLOBAL PORTS -----
input [0:0] SC1;
//----- GLOBAL PORTS -----
input [0:0] SR;
//----- GLOBAL PORTS -----
input [0:0] SE2;
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GPIN PORTS -----
input [0:93] gfpga_pad_pinput_extmode_A2F;
//----- GPIN PORTS -----
input [0:1] gfpga_pad_pinput_dchain_extmode_A2F;
//----- GPOUT PORTS -----
output [0:93] gfpga_pad_pinput_extmode_mode_o;
//----- GPOUT PORTS -----
output [0:95] gfpga_pad_poutput_F2A;
//----- GPOUT PORTS -----
output [0:11] gfpga_pad_mmffosc2cko_wrapper_C_O;
//----- GPOUT PORTS -----
output [0:1] gfpga_pad_pinput_dchain_extmode_mode_o;
//----- INPUT PORTS -----
input [0:7] ccff_head;
//----- OUTPUT PORTS -----
output [0:7] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:63] tile_0__0__undriven_cbx_0__chanx_left_in;
wire [0:63] tile_0__0__undriven_cbx_0__chanx_left_out;
wire [0:31] tile_0__0__undriven_cby_0__chany_bottom_in;
wire [0:31] tile_0__0__undriven_cby_0__chany_bottom_out;
wire [0:63] tile_0__1__undriven_cbx_0__chanx_left_in;
wire [0:63] tile_0__1__undriven_cbx_0__chanx_left_out;
wire [0:31] tile_0__2__undriven_cbx_0__chanx_left_in;
wire [0:63] tile_0__2__undriven_cbx_0__chanx_left_out;
wire [0:63] tile_0__3__undriven_cbx_0__chanx_left_in;
wire [0:63] tile_0__3__undriven_cbx_0__chanx_left_out;
wire [0:31] tile_0__4__undriven_cbx_0__chanx_left_in;
wire [0:31] tile_0__4__undriven_cbx_0__chanx_left_out;
wire [0:31] tile_0__5__undriven_cby_0__chany_top_in;
wire [0:31] tile_0__5__undriven_cby_0__chany_top_out;
wire [0:63] tile_0__EMPTY_id7__0_sb_0__chanx_right_out;
wire [0:63] tile_0__EMPTY_id7__0_sb_0__chany_top_out;
wire [0:63] tile_10__io_bottomL_bottom_id5__0_cbx_0__chanx_left_out;
wire [0:63] tile_10__io_bottomL_bottom_id5__0_sb_0__chanx_right_out;
wire [0:63] tile_10__io_bottomL_bottom_id5__0_sb_0__chany_top_out;
wire [0:63] tile_11__clb_id14__0_cbx_0__chanx_left_out;
wire [0:63] tile_11__clb_id14__0_cby_0__chany_bottom_out;
wire [0:63] tile_11__clb_id14__0_sb_0__chanx_right_out;
wire [0:63] tile_11__clb_id14__0_sb_0__chany_top_out;
wire [0:63] tile_11__clb_id14__1_cbx_0__chanx_left_out;
wire [0:63] tile_11__clb_id14__1_cby_0__chany_bottom_out;
wire [0:63] tile_11__clb_id14__1_sb_0__chanx_right_out;
wire [0:63] tile_11__clb_id14__1_sb_0__chany_top_out;
wire [0:63] tile_11__clb_id14__2_cbx_0__chanx_left_out;
wire [0:63] tile_11__clb_id14__2_cby_0__chany_bottom_out;
wire [0:63] tile_11__clb_id14__2_sb_0__chanx_right_out;
wire [0:63] tile_11__clb_id14__2_sb_0__chany_top_out;
wire [0:63] tile_12__clb_id15__0_cbx_0__chanx_left_out;
wire [0:63] tile_12__clb_id15__0_cby_0__chany_bottom_out;
wire [0:31] tile_12__clb_id15__0_sb_0__chanx_right_out;
wire [0:63] tile_12__clb_id15__0_sb_0__chany_top_out;
wire [0:63] tile_13__EMPTY_id4__0_cbx_0__chanx_left_out;
wire [0:63] tile_14__io_rightL_right_id3__0_cbx_0__chanx_left_out;
wire [0:63] tile_14__io_rightL_right_id3__1_cbx_0__chanx_left_out;
wire [0:63] tile_14__io_rightL_right_id3__2_cbx_0__chanx_left_out;
wire [0:31] tile_15__io_rightL_right_id2__0_cbx_0__chanx_left_out;
wire [0:63] tile_1__0__undriven_cby_0__chany_bottom_in;
wire [0:63] tile_1__0__undriven_cby_0__chany_bottom_out;
wire [0:63] tile_1__5__undriven_cby_0__chany_top_in;
wire [0:63] tile_1__5__undriven_cby_0__chany_top_out;
wire [0:63] tile_1__io_leftL_left_id8__0_cby_0__chany_bottom_out;
wire [0:63] tile_1__io_leftL_left_id8__0_sb_0__chanx_right_out;
wire [0:63] tile_1__io_leftL_left_id8__0_sb_0__chany_top_out;
wire [0:63] tile_2__0__undriven_cby_0__chany_bottom_in;
wire [0:63] tile_2__0__undriven_cby_0__chany_bottom_out;
wire [0:63] tile_2__5__undriven_cby_0__chany_top_in;
wire [0:63] tile_2__5__undriven_cby_0__chany_top_out;
wire [0:63] tile_2__io_leftL_left_id9__0_cby_0__chany_bottom_out;
wire [0:63] tile_2__io_leftL_left_id9__0_sb_0__chanx_right_out;
wire [0:63] tile_2__io_leftL_left_id9__0_sb_0__chany_top_out;
wire [0:63] tile_3__0__undriven_cbx_0__chanx_right_in;
wire [0:63] tile_3__0__undriven_cbx_0__chanx_right_out;
wire [0:63] tile_3__1__undriven_cbx_0__chanx_right_in;
wire [0:63] tile_3__1__undriven_cbx_0__chanx_right_out;
wire [0:63] tile_3__2__undriven_cbx_0__chanx_right_in;
wire [0:63] tile_3__2__undriven_cbx_0__chanx_right_out;
wire [0:63] tile_3__3__undriven_cbx_0__chanx_right_in;
wire [0:63] tile_3__3__undriven_cbx_0__chanx_right_out;
wire [0:31] tile_3__4__undriven_cbx_0__chanx_right_in;
wire [0:31] tile_3__4__undriven_cbx_0__chanx_right_out;
wire [0:63] tile_3__io_leftL_left_id10__0_cby_0__chany_bottom_out;
wire [0:63] tile_3__io_leftL_left_id10__0_sb_0__chanx_right_out;
wire [0:63] tile_3__io_leftL_left_id10__0_sb_0__chany_top_out;
wire [0:63] tile_4__io_leftL_left_id11__0_cby_0__chany_bottom_out;
wire [0:63] tile_4__io_leftL_left_id11__0_sb_0__chanx_right_out;
wire [0:31] tile_4__io_leftL_left_id11__0_sb_0__chany_top_out;
wire [0:31] tile_5__EMPTY_id0__0_cby_0__chany_bottom_out;
wire [0:63] tile_6__io_bottomL_bottom_id6__0_cbx_0__chanx_left_out;
wire [0:63] tile_6__io_bottomL_bottom_id6__0_sb_0__chanx_right_out;
wire [0:63] tile_6__io_bottomL_bottom_id6__0_sb_0__chany_top_out;
wire [0:63] tile_7__clb_id12__0_cbx_0__chanx_left_out;
wire [0:63] tile_7__clb_id12__0_cby_0__chany_bottom_out;
wire [0:63] tile_7__clb_id12__0_sb_0__chanx_right_out;
wire [0:63] tile_7__clb_id12__0_sb_0__chany_top_out;
wire [0:63] tile_7__clb_id12__1_cbx_0__chanx_left_out;
wire [0:63] tile_7__clb_id12__1_cby_0__chany_bottom_out;
wire [0:63] tile_7__clb_id12__1_sb_0__chanx_right_out;
wire [0:63] tile_7__clb_id12__1_sb_0__chany_top_out;
wire [0:63] tile_7__clb_id12__2_cbx_0__chanx_left_out;
wire [0:63] tile_7__clb_id12__2_cby_0__chany_bottom_out;
wire [0:63] tile_7__clb_id12__2_sb_0__chanx_right_out;
wire [0:63] tile_7__clb_id12__2_sb_0__chany_top_out;
wire [0:63] tile_8__clb_id13__0_cbx_0__chanx_left_out;
wire [0:63] tile_8__clb_id13__0_cby_0__chany_bottom_out;
wire [0:63] tile_8__clb_id13__0_sb_0__chanx_right_out;
wire [0:63] tile_8__clb_id13__0_sb_0__chany_top_out;
wire [0:63] tile_9__io_topL_top_id1__0_cby_0__chany_bottom_out;
wire [0:63] tile_9__io_topL_top_id1__1_cby_0__chany_bottom_out;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[0] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[1] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[2] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[3] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[4] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[5] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[6] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[7] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[8] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[9] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[10] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[11] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[12] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[13] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[14] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[15] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[16] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[17] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[18] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[19] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[20] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[21] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[22] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[23] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[24] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[25] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[26] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[27] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[28] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[29] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[30] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[31] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[32] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[33] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[34] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[35] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[36] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[37] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[38] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[39] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[40] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[41] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[42] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[43] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[44] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[45] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[46] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[47] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[48] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[49] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[50] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[51] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[52] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[53] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[54] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[55] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[56] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[57] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[58] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[59] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[60] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[61] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[62] = 1'b0;
	assign tile_0__0__undriven_cbx_0__chanx_left_in[63] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[0] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[1] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[2] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[3] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[4] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[5] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[6] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[7] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[8] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[9] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[10] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[11] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[12] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[13] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[14] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[15] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[16] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[17] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[18] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[19] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[20] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[21] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[22] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[23] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[24] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[25] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[26] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[27] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[28] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[29] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[30] = 1'b0;
	assign tile_0__0__undriven_cby_0__chany_bottom_in[31] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[0] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[1] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[2] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[3] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[4] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[5] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[6] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[7] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[8] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[9] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[10] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[11] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[12] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[13] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[14] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[15] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[16] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[17] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[18] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[19] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[20] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[21] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[22] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[23] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[24] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[25] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[26] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[27] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[28] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[29] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[30] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[31] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[32] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[33] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[34] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[35] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[36] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[37] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[38] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[39] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[40] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[41] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[42] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[43] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[44] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[45] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[46] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[47] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[48] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[49] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[50] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[51] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[52] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[53] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[54] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[55] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[56] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[57] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[58] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[59] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[60] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[61] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[62] = 1'b0;
	assign tile_0__1__undriven_cbx_0__chanx_left_in[63] = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[0] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[1] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[2] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[3] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[4] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[5] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[6] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[7] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[8] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[9] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[10] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[11] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[12] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[13] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[14] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[15] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[16] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[17] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[18] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[19] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[20] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[21] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[22] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[23] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[24] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[25] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[26] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[27] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[28] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[29] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[30] = 1'b0;
	assign tile_0__2__undriven_cbx_0__chanx_left_in[31] = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[0] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[1] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[2] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[3] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[4] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[5] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[6] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[7] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[8] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[9] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[10] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[11] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[12] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[13] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[14] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[15] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[16] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[17] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[18] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[19] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[20] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[21] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[22] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[23] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[24] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[25] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[26] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[27] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[28] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[29] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[30] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[31] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[32] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[33] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[34] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[35] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[36] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[37] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[38] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[39] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[40] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[41] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[42] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[43] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[44] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[45] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[46] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[47] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[48] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[49] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[50] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[51] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[52] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[53] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[54] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[55] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[56] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[57] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[58] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[59] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[60] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[61] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[62] = 1'b0;
	assign tile_0__3__undriven_cbx_0__chanx_left_in[63] = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[0] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[1] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[2] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[3] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[4] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[5] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[6] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[7] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[8] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[9] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[10] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[11] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[12] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[13] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[14] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[15] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[16] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[17] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[18] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[19] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[20] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[21] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[22] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[23] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[24] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[25] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[26] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[27] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[28] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[29] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[30] = 1'b0;
	assign tile_0__4__undriven_cbx_0__chanx_left_in[31] = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[0] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[1] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[2] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[3] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[4] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[5] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[6] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[7] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[8] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[9] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[10] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[11] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[12] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[13] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[14] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[15] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[16] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[17] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[18] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[19] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[20] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[21] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[22] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[23] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[24] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[25] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[26] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[27] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[28] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[29] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[30] = 1'b0;
	assign tile_0__5__undriven_cby_0__chany_top_in[31] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[0] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[1] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[2] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[3] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[4] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[5] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[6] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[7] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[8] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[9] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[10] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[11] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[12] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[13] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[14] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[15] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[16] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[17] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[18] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[19] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[20] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[21] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[22] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[23] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[24] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[25] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[26] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[27] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[28] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[29] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[30] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[31] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[32] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[33] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[34] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[35] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[36] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[37] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[38] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[39] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[40] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[41] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[42] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[43] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[44] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[45] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[46] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[47] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[48] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[49] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[50] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[51] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[52] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[53] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[54] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[55] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[56] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[57] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[58] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[59] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[60] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[61] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[62] = 1'b0;
	assign tile_1__0__undriven_cby_0__chany_bottom_in[63] = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_1__4__undriven_grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_ = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[0] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[1] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[2] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[3] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[4] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[5] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[6] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[7] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[8] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[9] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[10] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[11] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[12] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[13] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[14] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[15] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[16] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[17] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[18] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[19] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[20] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[21] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[22] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[23] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[24] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[25] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[26] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[27] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[28] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[29] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[30] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[31] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[32] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[33] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[34] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[35] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[36] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[37] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[38] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[39] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[40] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[41] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[42] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[43] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[44] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[45] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[46] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[47] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[48] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[49] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[50] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[51] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[52] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[53] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[54] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[55] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[56] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[57] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[58] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[59] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[60] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[61] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[62] = 1'b0;
	assign tile_1__5__undriven_cby_0__chany_top_in[63] = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[0] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[1] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[2] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[3] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[4] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[5] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[6] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[7] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[8] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[9] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[10] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[11] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[12] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[13] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[14] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[15] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[16] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[17] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[18] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[19] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[20] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[21] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[22] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[23] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[24] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[25] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[26] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[27] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[28] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[29] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[30] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[31] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[32] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[33] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[34] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[35] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[36] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[37] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[38] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[39] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[40] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[41] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[42] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[43] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[44] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[45] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[46] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[47] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[48] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[49] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[50] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[51] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[52] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[53] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[54] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[55] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[56] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[57] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[58] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[59] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[60] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[61] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[62] = 1'b0;
	assign tile_2__0__undriven_cby_0__chany_bottom_in[63] = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_2__4__undriven_grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_ = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[0] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[1] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[2] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[3] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[4] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[5] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[6] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[7] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[8] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[9] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[10] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[11] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[12] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[13] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[14] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[15] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[16] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[17] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[18] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[19] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[20] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[21] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[22] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[23] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[24] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[25] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[26] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[27] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[28] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[29] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[30] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[31] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[32] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[33] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[34] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[35] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[36] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[37] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[38] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[39] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[40] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[41] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[42] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[43] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[44] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[45] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[46] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[47] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[48] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[49] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[50] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[51] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[52] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[53] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[54] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[55] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[56] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[57] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[58] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[59] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[60] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[61] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[62] = 1'b0;
	assign tile_2__5__undriven_cby_0__chany_top_in[63] = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[0] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[1] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[2] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[3] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[4] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[5] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[6] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[7] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[8] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[9] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[10] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[11] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[12] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[13] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[14] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[15] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[16] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[17] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[18] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[19] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[20] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[21] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[22] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[23] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[24] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[25] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[26] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[27] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[28] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[29] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[30] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[31] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[32] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[33] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[34] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[35] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[36] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[37] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[38] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[39] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[40] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[41] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[42] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[43] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[44] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[45] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[46] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[47] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[48] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[49] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[50] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[51] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[52] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[53] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[54] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[55] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[56] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[57] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[58] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[59] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[60] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[61] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[62] = 1'b0;
	assign tile_3__0__undriven_cbx_0__chanx_right_in[63] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[0] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[1] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[2] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[3] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[4] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[5] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[6] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[7] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[8] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[9] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[10] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[11] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[12] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[13] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[14] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[15] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[16] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[17] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[18] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[19] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[20] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[21] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[22] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[23] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[24] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[25] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[26] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[27] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[28] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[29] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[30] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[31] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[32] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[33] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[34] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[35] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[36] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[37] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[38] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[39] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[40] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[41] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[42] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[43] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[44] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[45] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[46] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[47] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[48] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[49] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[50] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[51] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[52] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[53] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[54] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[55] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[56] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[57] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[58] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[59] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[60] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[61] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[62] = 1'b0;
	assign tile_3__1__undriven_cbx_0__chanx_right_in[63] = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[0] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[1] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[2] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[3] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[4] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[5] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[6] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[7] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[8] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[9] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[10] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[11] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[12] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[13] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[14] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[15] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[16] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[17] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[18] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[19] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[20] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[21] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[22] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[23] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[24] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[25] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[26] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[27] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[28] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[29] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[30] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[31] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[32] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[33] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[34] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[35] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[36] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[37] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[38] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[39] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[40] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[41] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[42] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[43] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[44] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[45] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[46] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[47] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[48] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[49] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[50] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[51] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[52] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[53] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[54] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[55] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[56] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[57] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[58] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[59] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[60] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[61] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[62] = 1'b0;
	assign tile_3__2__undriven_cbx_0__chanx_right_in[63] = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[0] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[1] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[2] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[3] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[4] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[5] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[6] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[7] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[8] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[9] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[10] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[11] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[12] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[13] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[14] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[15] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[16] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[17] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[18] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[19] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[20] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[21] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[22] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[23] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[24] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[25] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[26] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[27] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[28] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[29] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[30] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[31] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[32] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[33] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[34] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[35] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[36] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[37] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[38] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[39] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[40] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[41] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[42] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[43] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[44] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[45] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[46] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[47] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[48] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[49] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[50] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[51] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[52] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[53] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[54] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[55] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[56] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[57] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[58] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[59] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[60] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[61] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[62] = 1'b0;
	assign tile_3__3__undriven_cbx_0__chanx_right_in[63] = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[0] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[1] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[2] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[3] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[4] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[5] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[6] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[7] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[8] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[9] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[10] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[11] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[12] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[13] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[14] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[15] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[16] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[17] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[18] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[19] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[20] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[21] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[22] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[23] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[24] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[25] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[26] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[27] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[28] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[29] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[30] = 1'b0;
	assign tile_3__4__undriven_cbx_0__chanx_right_in[31] = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_ = 1'b0;
	assign tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_ = 1'b0;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	tile_5__EMPTY_id0_ tile_0__5_ (
		.cby_0__chany_bottom_in(tile_4__io_leftL_left_id11__0_sb_0__chany_top_out[0:31]),
		.cby_0__chany_top_in(tile_0__5__undriven_cby_0__chany_top_in[0:31]),
		.cby_0__chany_bottom_out(tile_5__EMPTY_id0__0_cby_0__chany_bottom_out[0:31]),
		.cby_0__chany_top_out(tile_0__5__undriven_cby_0__chany_top_out[0:31]));

	tile_9__io_topL_top_id1_ tile_1__5_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[7]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[0:7]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[0:7]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[0:7]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[0]),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_in_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cby_0__chany_bottom_in(tile_8__clb_id13__0_sb_0__chany_top_out[0:63]),
		.cby_0__chany_top_in(tile_1__5__undriven_cby_0__chany_top_in[0:63]),
		.ccff_head(tile_9__io_topL_top_id1__1_ccff_tail),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_out_0_(tile_1__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cby_0__chany_bottom_out(tile_9__io_topL_top_id1__0_cby_0__chany_bottom_out[0:63]),
		.cby_0__chany_top_out(tile_1__5__undriven_cby_0__chany_top_out[0:63]),
		.ccff_tail(ccff_tail[7]));

	tile_9__io_topL_top_id1_ tile_2__5_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[7]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[8:15]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[8:15]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[8:15]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[1]),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_in_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cby_0__chany_bottom_in(tile_12__clb_id15__0_sb_0__chany_top_out[0:63]),
		.cby_0__chany_top_in(tile_2__5__undriven_cby_0__chany_top_in[0:63]),
		.ccff_head(tile_15__io_rightL_right_id2__0_ccff_tail),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_out_0_(tile_2__5__undriven_grid_io_topL_top_bottom_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cby_0__chany_bottom_out(tile_9__io_topL_top_id1__1_cby_0__chany_bottom_out[0:63]),
		.cby_0__chany_top_out(tile_2__5__undriven_cby_0__chany_top_out[0:63]),
		.ccff_tail(tile_9__io_topL_top_id1__1_ccff_tail));

	tile_15__io_rightL_right_id2_ tile_3__4_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[7]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[16:23]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[16:23]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[16:23]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[2]),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.cbx_0__chanx_left_in(tile_12__clb_id15__0_sb_0__chanx_right_out[0:31]),
		.cbx_0__chanx_right_in(tile_3__4__undriven_cbx_0__chanx_right_in[0:31]),
		.ccff_head(tile_12__clb_id15__0_ccff_tail),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_(tile_3__4__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_15__io_rightL_right_id2__0_cbx_0__chanx_left_out[0:31]),
		.cbx_0__chanx_right_out(tile_3__4__undriven_cbx_0__chanx_right_out[0:31]),
		.ccff_tail(tile_15__io_rightL_right_id2__0_ccff_tail));

	tile_14__io_rightL_right_id3_ tile_3__3_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[5]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[24:31]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[24:31]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[24:31]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[3]),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.cbx_0__chanx_left_in(tile_11__clb_id14__2_sb_0__chanx_right_out[0:63]),
		.cbx_0__chanx_right_in(tile_3__3__undriven_cbx_0__chanx_right_in[0:63]),
		.ccff_head(tile_14__io_rightL_right_id3__1_ccff_tail),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_(tile_3__3__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_14__io_rightL_right_id3__0_cbx_0__chanx_left_out[0:63]),
		.cbx_0__chanx_right_out(tile_3__3__undriven_cbx_0__chanx_right_out[0:63]),
		.ccff_tail(ccff_tail[5]));

	tile_14__io_rightL_right_id3_ tile_3__2_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[5]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[32:39]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[32:39]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[32:39]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[4]),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.cbx_0__chanx_left_in(tile_11__clb_id14__1_sb_0__chanx_right_out[0:63]),
		.cbx_0__chanx_right_in(tile_3__2__undriven_cbx_0__chanx_right_in[0:63]),
		.ccff_head(ccff_head[5]),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_(tile_3__2__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_14__io_rightL_right_id3__1_cbx_0__chanx_left_out[0:63]),
		.cbx_0__chanx_right_out(tile_3__2__undriven_cbx_0__chanx_right_out[0:63]),
		.ccff_tail(tile_14__io_rightL_right_id3__1_ccff_tail));

	tile_14__io_rightL_right_id3_ tile_3__1_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[1]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[40:47]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[40:47]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[40:47]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[5]),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_in_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.cbx_0__chanx_left_in(tile_11__clb_id14__0_sb_0__chanx_right_out[0:63]),
		.cbx_0__chanx_right_in(tile_3__1__undriven_cbx_0__chanx_right_in[0:63]),
		.ccff_head(tile_10__io_bottomL_bottom_id5__0_ccff_tail),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_(tile_3__1__undriven_grid_io_rightL_right_left_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_14__io_rightL_right_id3__2_cbx_0__chanx_left_out[0:63]),
		.cbx_0__chanx_right_out(tile_3__1__undriven_cbx_0__chanx_right_out[0:63]),
		.ccff_tail(ccff_tail[1]));

	tile_13__EMPTY_id4_ tile_3__0_ (
		.cbx_0__chanx_left_in(tile_10__io_bottomL_bottom_id5__0_sb_0__chanx_right_out[0:63]),
		.cbx_0__chanx_right_in(tile_3__0__undriven_cbx_0__chanx_right_in[0:63]),
		.cbx_0__chanx_left_out(tile_13__EMPTY_id4__0_cbx_0__chanx_left_out[0:63]),
		.cbx_0__chanx_right_out(tile_3__0__undriven_cbx_0__chanx_right_out[0:63]));

	tile_10__io_bottomL_bottom_id5_ tile_2__0_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[1]),
		.gfpga_pad_pinput_dchain_extmode_A2F(gfpga_pad_pinput_dchain_extmode_A2F[0]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[48:54]),
		.gfpga_pad_pinput_dchain_extmode_mode_o(gfpga_pad_pinput_dchain_extmode_mode_o[0]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[48:54]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[48:55]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[6]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_11__clb_id14__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_13__EMPTY_id4__0_cbx_0__chanx_left_out[0:63]),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_in_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cbx_0__chanx_left_in(tile_6__io_bottomL_bottom_id6__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_2__0__undriven_cby_0__chany_bottom_in[0:63]),
		.ccff_head(ccff_head[1]),
		.sb_0__chany_top_out(tile_10__io_bottomL_bottom_id5__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_10__io_bottomL_bottom_id5__0_sb_0__chanx_right_out[0:63]),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_out_0_(tile_2__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_10__io_bottomL_bottom_id5__0_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_2__0__undriven_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_10__io_bottomL_bottom_id5__0_ccff_tail));

	tile_6__io_bottomL_bottom_id6_ tile_1__0_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_pinput_dchain_extmode_A2F(gfpga_pad_pinput_dchain_extmode_A2F[1]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[55:61]),
		.gfpga_pad_pinput_dchain_extmode_mode_o(gfpga_pad_pinput_dchain_extmode_mode_o[1]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[55:61]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[56:63]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[7]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_10__io_bottomL_bottom_id5__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_7__clb_id12__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_10__io_bottomL_bottom_id5__0_cbx_0__chanx_left_out[0:63]),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_in_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cbx_0__chanx_left_in(tile_0__EMPTY_id7__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_1__0__undriven_cby_0__chany_bottom_in[0:63]),
		.ccff_head(tile_0__EMPTY_id7__0_ccff_tail),
		.sb_0__chany_top_out(tile_6__io_bottomL_bottom_id6__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_6__io_bottomL_bottom_id6__0_sb_0__chanx_right_out[0:63]),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_out_0_(tile_1__0__undriven_grid_io_bottomL_bottom_top_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_6__io_bottomL_bottom_id6__0_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_1__0__undriven_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(ccff_tail[0]));

	tile_0__EMPTY_id7_ tile_0__0_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[0]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_6__io_bottomL_bottom_id6__0_grid_io_bottomL_bottom_top_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_1__io_leftL_left_id8__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_6__io_bottomL_bottom_id6__0_cbx_0__chanx_left_out[0:63]),
		.cbx_0__chanx_left_in(tile_0__0__undriven_cbx_0__chanx_left_in[0:63]),
		.cby_0__chany_bottom_in(tile_0__0__undriven_cby_0__chany_bottom_in[0:31]),
		.ccff_head(ccff_head[0]),
		.sb_0__chany_top_out(tile_0__EMPTY_id7__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_0__EMPTY_id7__0_sb_0__chanx_right_out[0:63]),
		.cbx_0__chanx_left_out(tile_0__0__undriven_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_0__0__undriven_cby_0__chany_bottom_out[0:31]),
		.ccff_tail(tile_0__EMPTY_id7__0_ccff_tail));

	tile_1__io_leftL_left_id8_ tile_0__1_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[3]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[62:69]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[62:69]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[64:71]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[8]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_4__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_5__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_6__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_7__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_8__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_9__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_10__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_11__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_12__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_13__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_14__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_15__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_16__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_17__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_18__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_19__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__chany_top_in(tile_2__io_leftL_left_id9__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_7__clb_id12__0_cbx_0__chanx_left_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cbx_0__chanx_left_in(tile_0__1__undriven_cbx_0__chanx_left_in[0:63]),
		.cby_0__chany_bottom_in(tile_0__EMPTY_id7__0_sb_0__chany_top_out[0:63]),
		.ccff_head(ccff_head[3]),
		.sb_0__chany_top_out(tile_1__io_leftL_left_id8__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_1__io_leftL_left_id8__0_sb_0__chanx_right_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_1__io_leftL_left_id8__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_(tile_0__1__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_0__1__undriven_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_1__io_leftL_left_id8__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_1__io_leftL_left_id8__0_ccff_tail));

	tile_2__io_leftL_left_id9_ tile_0__2_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[3]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[70:77]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[70:77]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[72:79]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[9]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_4__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_5__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_6__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_7__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_8__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_9__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_10__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_11__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_12__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_13__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_14__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_15__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_16__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_17__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_18__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_19__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_4__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_5__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_6__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_7__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_8__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_9__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_10__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_11__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_12__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_13__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_14__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_15__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_16__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_17__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_18__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_19__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.sb_0__chany_top_in(tile_3__io_leftL_left_id10__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_7__clb_id12__1_cbx_0__chanx_left_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cbx_0__chanx_left_in({tile_0__2__undriven_cbx_0__chanx_left_in[0:31], clk[0:7], reset[0:23]}),
		.cby_0__chany_bottom_in(tile_1__io_leftL_left_id8__0_sb_0__chany_top_out[0:63]),
		.ccff_head(tile_1__io_leftL_left_id8__0_ccff_tail),
		.sb_0__chany_top_out(tile_2__io_leftL_left_id9__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_2__io_leftL_left_id9__0_sb_0__chanx_right_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_2__io_leftL_left_id9__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_(tile_0__2__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_0__2__undriven_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_2__io_leftL_left_id9__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(ccff_tail[3]));

	tile_3__io_leftL_left_id10_ tile_0__3_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[7]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[78:85]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[78:85]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[80:87]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[10]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_4__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_5__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_6__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_7__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_8__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_9__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_10__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_11__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_12__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_13__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_14__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_15__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_16__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_17__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_18__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_19__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.sb_0__chany_top_in(tile_4__io_leftL_left_id11__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_7__clb_id12__2_cbx_0__chanx_left_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cbx_0__chanx_left_in(tile_0__3__undriven_cbx_0__chanx_left_in[0:63]),
		.cby_0__chany_bottom_in(tile_2__io_leftL_left_id9__0_sb_0__chany_top_out[0:63]),
		.ccff_head(ccff_head[7]),
		.sb_0__chany_top_out(tile_3__io_leftL_left_id10__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_3__io_leftL_left_id10__0_sb_0__chanx_right_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_3__io_leftL_left_id10__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_(tile_0__3__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_0__3__undriven_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_3__io_leftL_left_id10__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_3__io_leftL_left_id10__0_ccff_tail));

	tile_4__io_leftL_left_id11_ tile_0__4_ (
		.SE0(SE0),
		.SE1(SE1),
		.SC0(SC0),
		.SC1(SC1),
		.SR(SR),
		.SE2(SE2),
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[7]),
		.gfpga_pad_pinput_extmode_A2F(gfpga_pad_pinput_extmode_A2F[86:93]),
		.gfpga_pad_pinput_extmode_mode_o(gfpga_pad_pinput_extmode_mode_o[86:93]),
		.gfpga_pad_poutput_F2A(gfpga_pad_poutput_F2A[88:95]),
		.gfpga_pad_mmffosc2cko_wrapper_C_O(gfpga_pad_mmffosc2cko_wrapper_C_O[11]),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__chany_top_in(tile_5__EMPTY_id0__0_cby_0__chany_bottom_out[0:31]),
		.sb_0__chanx_right_in(tile_8__clb_id13__0_cbx_0__chanx_left_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_in_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_in_0_),
		.cbx_0__chanx_left_in(tile_0__4__undriven_cbx_0__chanx_left_in[0:31]),
		.cby_0__chany_bottom_in(tile_3__io_leftL_left_id10__0_sb_0__chany_top_out[0:63]),
		.ccff_head(tile_3__io_leftL_left_id10__0_ccff_tail),
		.sb_0__chany_top_out(tile_4__io_leftL_left_id11__0_sb_0__chany_top_out[0:31]),
		.sb_0__chanx_right_out(tile_4__io_leftL_left_id11__0_sb_0__chanx_right_out[0:63]),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_0__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_1__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_2__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_3__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_4__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_5__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_6__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_4__io_leftL_left_id11__0_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_7__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_8__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_9__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_10__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_11__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_12__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_13__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_14__pin_sc_out_0_),
		.grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_(tile_0__4__undriven_grid_io_leftL_left_right_width_0_height_0_subtile_15__pin_sc_out_0_),
		.cbx_0__chanx_left_out(tile_0__4__undriven_cbx_0__chanx_left_out[0:31]),
		.cby_0__chany_bottom_out(tile_4__io_leftL_left_id11__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_4__io_leftL_left_id11__0_ccff_tail));

	tile_7__clb_id12_ tile_1__1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[2]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__chany_top_in(tile_7__clb_id12__1_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_11__clb_id14__0_cbx_0__chanx_left_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_0_out),
		.cbx_0__chanx_left_in(tile_1__io_leftL_left_id8__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_6__io_bottomL_bottom_id6__0_sb_0__chany_top_out[0:63]),
		.ccff_head(tile_11__clb_id14__0_ccff_tail),
		.sb_0__chany_top_out(tile_7__clb_id12__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_7__clb_id12__0_sb_0__chanx_right_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_7__clb_id12__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_7__clb_id12__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_1__1__undriven_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_1__1__undriven_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_7__clb_id12__0_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_7__clb_id12__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(ccff_tail[2]));

	tile_7__clb_id12_ tile_1__2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[4]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__chany_top_in(tile_7__clb_id12__2_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_11__clb_id14__1_cbx_0__chanx_left_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_1_out),
		.cbx_0__chanx_left_in(tile_2__io_leftL_left_id9__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_7__clb_id12__0_sb_0__chany_top_out[0:63]),
		.ccff_head(ccff_head[4]),
		.sb_0__chany_top_out(tile_7__clb_id12__1_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_7__clb_id12__1_sb_0__chanx_right_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_7__clb_id12__1_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_7__clb_id12__1_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_7__clb_id12__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_7__clb_id12__1_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_7__clb_id12__1_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_7__clb_id12__1_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_7__clb_id12__1_ccff_tail));

	tile_7__clb_id12_ tile_1__3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[6]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__chany_top_in(tile_8__clb_id13__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_11__clb_id14__2_cbx_0__chanx_left_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_2_out),
		.cbx_0__chanx_left_in(tile_3__io_leftL_left_id10__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_7__clb_id12__1_sb_0__chany_top_out[0:63]),
		.ccff_head(tile_11__clb_id14__2_ccff_tail),
		.sb_0__chany_top_out(tile_7__clb_id12__2_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_7__clb_id12__2_sb_0__chanx_right_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_7__clb_id12__2_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_7__clb_id12__2_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_7__clb_id12__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_7__clb_id12__2_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_7__clb_id12__2_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_7__clb_id12__2_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(ccff_tail[6]));

	tile_8__clb_id13_ tile_1__4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[7]),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__right_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.sb_0__right_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_9__io_topL_top_id1__0_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_9__io_topL_top_id1__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_12__clb_id15__0_cbx_0__chanx_left_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(tile_1__4__undriven_grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_),
		.cbx_0__chanx_left_in(tile_4__io_leftL_left_id11__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_7__clb_id12__2_sb_0__chany_top_out[0:63]),
		.ccff_head(tile_4__io_leftL_left_id11__0_ccff_tail),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_8__clb_id13__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.sb_0__chany_top_out(tile_8__clb_id13__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_8__clb_id13__0_sb_0__chanx_right_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_8__clb_id13__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_8__clb_id13__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_8__clb_id13__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_1__4__undriven_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_8__clb_id13__0_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_8__clb_id13__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_8__clb_id13__0_ccff_tail));

	tile_11__clb_id14_ tile_2__1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[2]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__2_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_11__clb_id14__1_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_14__io_rightL_right_id3__2_cbx_0__chanx_left_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_3_out),
		.cbx_0__chanx_left_in(tile_7__clb_id12__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_10__io_bottomL_bottom_id5__0_sb_0__chany_top_out[0:63]),
		.ccff_head(ccff_head[2]),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_(tile_11__clb_id14__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.sb_0__chany_top_out(tile_11__clb_id14__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_11__clb_id14__0_sb_0__chanx_right_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_11__clb_id14__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_11__clb_id14__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_2__1__undriven_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_2__1__undriven_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_11__clb_id14__0_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_11__clb_id14__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_11__clb_id14__0_ccff_tail));

	tile_11__clb_id14_ tile_2__2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[4]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__1_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_11__clb_id14__2_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_14__io_rightL_right_id3__1_cbx_0__chanx_left_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_4_out),
		.cbx_0__chanx_left_in(tile_7__clb_id12__1_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_11__clb_id14__0_sb_0__chany_top_out[0:63]),
		.ccff_head(tile_7__clb_id12__1_ccff_tail),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_(tile_11__clb_id14__1_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.sb_0__chany_top_out(tile_11__clb_id14__1_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_11__clb_id14__1_sb_0__chanx_right_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_11__clb_id14__1_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_11__clb_id14__1_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_11__clb_id14__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_2__2__undriven_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_11__clb_id14__1_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_11__clb_id14__1_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(ccff_tail[4]));

	tile_11__clb_id14_ tile_2__3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[6]),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_2_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_4_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_6_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_7_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.sb_0__top_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__top_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_14__io_rightL_right_id3__0_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_12__clb_id15__0_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_14__io_rightL_right_id3__0_cbx_0__chanx_left_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_5_out),
		.cbx_0__chanx_left_in(tile_7__clb_id12__2_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_11__clb_id14__1_sb_0__chany_top_out[0:63]),
		.ccff_head(ccff_head[6]),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_(tile_11__clb_id14__2_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.sb_0__chany_top_out(tile_11__clb_id14__2_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_11__clb_id14__2_sb_0__chanx_right_out[0:63]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_11__clb_id14__2_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_11__clb_id14__2_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_11__clb_id14__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_2__3__undriven_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_11__clb_id14__2_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_11__clb_id14__2_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_11__clb_id14__2_ccff_tail));

	tile_12__clb_id15_ tile_2__4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk[7]),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_15__io_rightL_right_id2__0_grid_io_rightL_right_left_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_),
		.sb_0__left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_(tile_9__io_topL_top_id1__1_grid_io_topL_top_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_),
		.sb_0__chany_top_in(tile_9__io_topL_top_id1__1_cby_0__chany_bottom_out[0:63]),
		.sb_0__chanx_right_in(tile_15__io_rightL_right_id2__0_cbx_0__chanx_left_out[0:31]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_(tile_2__4__undriven_grid_clb_top_width_0_height_0_subtile_0__pin_cin_0_),
		.cbx_0__chanx_left_in(tile_8__clb_id13__0_sb_0__chanx_right_out[0:63]),
		.cby_0__chany_bottom_in(tile_11__clb_id14__2_sb_0__chany_top_out[0:63]),
		.ccff_head(tile_8__clb_id13__0_ccff_tail),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.cbx_0__top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_12__clb_id15__0_cbx_0__top_grid_bottom_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_0__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_1__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_2__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_3__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_4__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_5__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_6__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_7__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_8__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_9__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_10__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_11__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_12__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_13__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_14__pin_clk_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_f2a_i_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_reset_0_),
		.cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_(tile_12__clb_id15__0_cby_0__right_grid_left_width_0_height_0_subtile_15__pin_clk_0_),
		.sb_0__chany_top_out(tile_12__clb_id15__0_sb_0__chany_top_out[0:63]),
		.sb_0__chanx_right_out(tile_12__clb_id15__0_sb_0__chanx_right_out[0:31]),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_12_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_12_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_13_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_13_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_14_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_14_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_15_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_15_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_16_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_16_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_17_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_17_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_18_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_18_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_19_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_19_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_20_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_20_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_21_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_21_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_22_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_22_),
		.grid_clb_top_width_0_height_0_subtile_0__pin_O_23_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_0__pin_O_23_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_1__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_1__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_2__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_2__pin_zero_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_3__pin_match1_o_0_),
		.grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_(tile_12__clb_id15__0_grid_clb_top_width_0_height_0_subtile_3__pin_zero_o_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_0_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_1_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_1_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_2_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_2_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_3_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_3_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_4_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_4_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_5_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_5_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_6_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_6_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_7_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_7_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_8_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_8_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_9_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_9_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_10_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_10_),
		.grid_clb_right_width_0_height_0_subtile_0__pin_O_11_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_0__pin_O_11_),
		.grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_1__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_2__pin_match0_o_0_),
		.grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_(tile_12__clb_id15__0_grid_clb_right_width_0_height_0_subtile_3__pin_match0_o_0_),
		.grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_(tile_12__clb_id15__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.grid_clb_left_width_0_height_0_subtile_4__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_4__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_5__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_5__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_6__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_6__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_7__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_7__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_8__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_8__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_9__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_9__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_10__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_10__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_11__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_11__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_12__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_12__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_13__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_13__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_14__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_14__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_15__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_15__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_16__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_16__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_17__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_17__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_18__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_18__pin_out_0_),
		.grid_clb_left_width_0_height_0_subtile_19__pin_out_0_(tile_2__4__undriven_grid_clb_left_width_0_height_0_subtile_19__pin_out_0_),
		.cbx_0__chanx_left_out(tile_12__clb_id15__0_cbx_0__chanx_left_out[0:63]),
		.cby_0__chany_bottom_out(tile_12__clb_id15__0_cby_0__chany_bottom_out[0:63]),
		.ccff_tail(tile_12__clb_id15__0_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(tile_7__clb_id12__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(tile_7__clb_id12__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(tile_8__clb_id13__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(tile_11__clb_id14__1_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(tile_11__clb_id14__2_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(tile_12__clb_id15__0_grid_clb_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_5_out));

endmodule
// ----- END Verilog module for fpga_core -----




