//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[2][4]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for sb_12_ -----
module sb_12_(config_enable,
              prog_reset,
              prog_clk,
              chany_top_in,
              chanx_right_in,
              chany_bottom_in,
              bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_,
              bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_,
              bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_,
              bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_,
              bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_,
              bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_,
              bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_,
              bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_,
              bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_,
              bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_,
              bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_,
              bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_,
              chanx_left_in,
              left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_,
              left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_,
              left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_,
              left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_,
              left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_,
              left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_,
              left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_,
              left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_,
              left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_,
              left_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_,
              left_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_,
              left_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_,
              left_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_,
              left_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_,
              left_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_,
              ccff_head,
              chany_top_out,
              chanx_right_out,
              chany_bottom_out,
              chanx_left_out,
              ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:63] chany_top_in;
//----- INPUT PORTS -----
input [0:31] chanx_right_in;
//----- INPUT PORTS -----
input [0:63] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_;
//----- INPUT PORTS -----
input [0:63] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:63] chany_top_out;
//----- OUTPUT PORTS -----
output [0:31] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:63] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:63] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] clk_mux_size3_0_sram;
wire [0:1] clk_mux_size3_0_sram_inv;
wire [0:1] clk_mux_size3_10_sram;
wire [0:1] clk_mux_size3_10_sram_inv;
wire [0:1] clk_mux_size3_11_sram;
wire [0:1] clk_mux_size3_11_sram_inv;
wire [0:1] clk_mux_size3_12_sram;
wire [0:1] clk_mux_size3_12_sram_inv;
wire [0:1] clk_mux_size3_13_sram;
wire [0:1] clk_mux_size3_13_sram_inv;
wire [0:1] clk_mux_size3_14_sram;
wire [0:1] clk_mux_size3_14_sram_inv;
wire [0:1] clk_mux_size3_15_sram;
wire [0:1] clk_mux_size3_15_sram_inv;
wire [0:1] clk_mux_size3_16_sram;
wire [0:1] clk_mux_size3_16_sram_inv;
wire [0:1] clk_mux_size3_17_sram;
wire [0:1] clk_mux_size3_17_sram_inv;
wire [0:1] clk_mux_size3_18_sram;
wire [0:1] clk_mux_size3_18_sram_inv;
wire [0:1] clk_mux_size3_19_sram;
wire [0:1] clk_mux_size3_19_sram_inv;
wire [0:1] clk_mux_size3_1_sram;
wire [0:1] clk_mux_size3_1_sram_inv;
wire [0:1] clk_mux_size3_20_sram;
wire [0:1] clk_mux_size3_20_sram_inv;
wire [0:1] clk_mux_size3_21_sram;
wire [0:1] clk_mux_size3_21_sram_inv;
wire [0:1] clk_mux_size3_22_sram;
wire [0:1] clk_mux_size3_22_sram_inv;
wire [0:1] clk_mux_size3_23_sram;
wire [0:1] clk_mux_size3_23_sram_inv;
wire [0:1] clk_mux_size3_24_sram;
wire [0:1] clk_mux_size3_24_sram_inv;
wire [0:1] clk_mux_size3_25_sram;
wire [0:1] clk_mux_size3_25_sram_inv;
wire [0:1] clk_mux_size3_26_sram;
wire [0:1] clk_mux_size3_26_sram_inv;
wire [0:1] clk_mux_size3_27_sram;
wire [0:1] clk_mux_size3_27_sram_inv;
wire [0:1] clk_mux_size3_28_sram;
wire [0:1] clk_mux_size3_28_sram_inv;
wire [0:1] clk_mux_size3_29_sram;
wire [0:1] clk_mux_size3_29_sram_inv;
wire [0:1] clk_mux_size3_2_sram;
wire [0:1] clk_mux_size3_2_sram_inv;
wire [0:1] clk_mux_size3_30_sram;
wire [0:1] clk_mux_size3_30_sram_inv;
wire [0:1] clk_mux_size3_31_sram;
wire [0:1] clk_mux_size3_31_sram_inv;
wire [0:1] clk_mux_size3_32_sram;
wire [0:1] clk_mux_size3_32_sram_inv;
wire [0:1] clk_mux_size3_33_sram;
wire [0:1] clk_mux_size3_33_sram_inv;
wire [0:1] clk_mux_size3_34_sram;
wire [0:1] clk_mux_size3_34_sram_inv;
wire [0:1] clk_mux_size3_35_sram;
wire [0:1] clk_mux_size3_35_sram_inv;
wire [0:1] clk_mux_size3_36_sram;
wire [0:1] clk_mux_size3_36_sram_inv;
wire [0:1] clk_mux_size3_37_sram;
wire [0:1] clk_mux_size3_37_sram_inv;
wire [0:1] clk_mux_size3_38_sram;
wire [0:1] clk_mux_size3_38_sram_inv;
wire [0:1] clk_mux_size3_39_sram;
wire [0:1] clk_mux_size3_39_sram_inv;
wire [0:1] clk_mux_size3_3_sram;
wire [0:1] clk_mux_size3_3_sram_inv;
wire [0:1] clk_mux_size3_40_sram;
wire [0:1] clk_mux_size3_40_sram_inv;
wire [0:1] clk_mux_size3_41_sram;
wire [0:1] clk_mux_size3_41_sram_inv;
wire [0:1] clk_mux_size3_42_sram;
wire [0:1] clk_mux_size3_42_sram_inv;
wire [0:1] clk_mux_size3_43_sram;
wire [0:1] clk_mux_size3_43_sram_inv;
wire [0:1] clk_mux_size3_44_sram;
wire [0:1] clk_mux_size3_44_sram_inv;
wire [0:1] clk_mux_size3_45_sram;
wire [0:1] clk_mux_size3_45_sram_inv;
wire [0:1] clk_mux_size3_46_sram;
wire [0:1] clk_mux_size3_46_sram_inv;
wire [0:1] clk_mux_size3_47_sram;
wire [0:1] clk_mux_size3_47_sram_inv;
wire [0:1] clk_mux_size3_48_sram;
wire [0:1] clk_mux_size3_48_sram_inv;
wire [0:1] clk_mux_size3_49_sram;
wire [0:1] clk_mux_size3_49_sram_inv;
wire [0:1] clk_mux_size3_4_sram;
wire [0:1] clk_mux_size3_4_sram_inv;
wire [0:1] clk_mux_size3_50_sram;
wire [0:1] clk_mux_size3_50_sram_inv;
wire [0:1] clk_mux_size3_51_sram;
wire [0:1] clk_mux_size3_51_sram_inv;
wire [0:1] clk_mux_size3_52_sram;
wire [0:1] clk_mux_size3_52_sram_inv;
wire [0:1] clk_mux_size3_53_sram;
wire [0:1] clk_mux_size3_53_sram_inv;
wire [0:1] clk_mux_size3_54_sram;
wire [0:1] clk_mux_size3_54_sram_inv;
wire [0:1] clk_mux_size3_55_sram;
wire [0:1] clk_mux_size3_55_sram_inv;
wire [0:1] clk_mux_size3_56_sram;
wire [0:1] clk_mux_size3_56_sram_inv;
wire [0:1] clk_mux_size3_57_sram;
wire [0:1] clk_mux_size3_57_sram_inv;
wire [0:1] clk_mux_size3_58_sram;
wire [0:1] clk_mux_size3_58_sram_inv;
wire [0:1] clk_mux_size3_59_sram;
wire [0:1] clk_mux_size3_59_sram_inv;
wire [0:1] clk_mux_size3_5_sram;
wire [0:1] clk_mux_size3_5_sram_inv;
wire [0:1] clk_mux_size3_60_sram;
wire [0:1] clk_mux_size3_60_sram_inv;
wire [0:1] clk_mux_size3_61_sram;
wire [0:1] clk_mux_size3_61_sram_inv;
wire [0:1] clk_mux_size3_62_sram;
wire [0:1] clk_mux_size3_62_sram_inv;
wire [0:1] clk_mux_size3_63_sram;
wire [0:1] clk_mux_size3_63_sram_inv;
wire [0:1] clk_mux_size3_6_sram;
wire [0:1] clk_mux_size3_6_sram_inv;
wire [0:1] clk_mux_size3_7_sram;
wire [0:1] clk_mux_size3_7_sram_inv;
wire [0:1] clk_mux_size3_8_sram;
wire [0:1] clk_mux_size3_8_sram_inv;
wire [0:1] clk_mux_size3_9_sram;
wire [0:1] clk_mux_size3_9_sram_inv;
wire [0:314] sb_12__config_group_mem_size315_0_mem_out;
wire [0:314] sb_12__config_group_mem_size315_0_mem_outb;
wire [0:3] sb_mux_size10_0_sram;
wire [0:3] sb_mux_size10_0_sram_inv;
wire [0:3] sb_mux_size10_1_sram;
wire [0:3] sb_mux_size10_1_sram_inv;
wire [0:3] sb_mux_size11_0_sram;
wire [0:3] sb_mux_size11_0_sram_inv;
wire [0:3] sb_mux_size11_1_sram;
wire [0:3] sb_mux_size11_1_sram_inv;
wire [0:3] sb_mux_size11_2_sram;
wire [0:3] sb_mux_size11_2_sram_inv;
wire [0:3] sb_mux_size11_3_sram;
wire [0:3] sb_mux_size11_3_sram_inv;
wire [0:1] sb_mux_size2_0_sram;
wire [0:1] sb_mux_size2_0_sram_inv;
wire [0:1] sb_mux_size2_10_sram;
wire [0:1] sb_mux_size2_10_sram_inv;
wire [0:1] sb_mux_size2_11_sram;
wire [0:1] sb_mux_size2_11_sram_inv;
wire [0:1] sb_mux_size2_12_sram;
wire [0:1] sb_mux_size2_12_sram_inv;
wire [0:1] sb_mux_size2_1_sram;
wire [0:1] sb_mux_size2_1_sram_inv;
wire [0:1] sb_mux_size2_2_sram;
wire [0:1] sb_mux_size2_2_sram_inv;
wire [0:1] sb_mux_size2_3_sram;
wire [0:1] sb_mux_size2_3_sram_inv;
wire [0:1] sb_mux_size2_4_sram;
wire [0:1] sb_mux_size2_4_sram_inv;
wire [0:1] sb_mux_size2_5_sram;
wire [0:1] sb_mux_size2_5_sram_inv;
wire [0:1] sb_mux_size2_6_sram;
wire [0:1] sb_mux_size2_6_sram_inv;
wire [0:1] sb_mux_size2_7_sram;
wire [0:1] sb_mux_size2_7_sram_inv;
wire [0:1] sb_mux_size2_8_sram;
wire [0:1] sb_mux_size2_8_sram_inv;
wire [0:1] sb_mux_size2_9_sram;
wire [0:1] sb_mux_size2_9_sram_inv;
wire [0:2] sb_mux_size4_0_sram;
wire [0:2] sb_mux_size4_0_sram_inv;
wire [0:2] sb_mux_size4_1_sram;
wire [0:2] sb_mux_size4_1_sram_inv;
wire [0:2] sb_mux_size4_2_sram;
wire [0:2] sb_mux_size4_2_sram_inv;
wire [0:2] sb_mux_size5_0_sram;
wire [0:2] sb_mux_size5_0_sram_inv;
wire [0:2] sb_mux_size5_1_sram;
wire [0:2] sb_mux_size5_1_sram_inv;
wire [0:2] sb_mux_size5_2_sram;
wire [0:2] sb_mux_size5_2_sram_inv;
wire [0:2] sb_mux_size6_0_sram;
wire [0:2] sb_mux_size6_0_sram_inv;
wire [0:2] sb_mux_size6_1_sram;
wire [0:2] sb_mux_size6_1_sram_inv;
wire [0:2] sb_mux_size7_0_sram;
wire [0:2] sb_mux_size7_0_sram_inv;
wire [0:2] sb_mux_size7_10_sram;
wire [0:2] sb_mux_size7_10_sram_inv;
wire [0:2] sb_mux_size7_11_sram;
wire [0:2] sb_mux_size7_11_sram_inv;
wire [0:2] sb_mux_size7_12_sram;
wire [0:2] sb_mux_size7_12_sram_inv;
wire [0:2] sb_mux_size7_13_sram;
wire [0:2] sb_mux_size7_13_sram_inv;
wire [0:2] sb_mux_size7_14_sram;
wire [0:2] sb_mux_size7_14_sram_inv;
wire [0:2] sb_mux_size7_1_sram;
wire [0:2] sb_mux_size7_1_sram_inv;
wire [0:2] sb_mux_size7_2_sram;
wire [0:2] sb_mux_size7_2_sram_inv;
wire [0:2] sb_mux_size7_3_sram;
wire [0:2] sb_mux_size7_3_sram_inv;
wire [0:2] sb_mux_size7_4_sram;
wire [0:2] sb_mux_size7_4_sram_inv;
wire [0:2] sb_mux_size7_5_sram;
wire [0:2] sb_mux_size7_5_sram_inv;
wire [0:2] sb_mux_size7_6_sram;
wire [0:2] sb_mux_size7_6_sram_inv;
wire [0:2] sb_mux_size7_7_sram;
wire [0:2] sb_mux_size7_7_sram_inv;
wire [0:2] sb_mux_size7_8_sram;
wire [0:2] sb_mux_size7_8_sram_inv;
wire [0:2] sb_mux_size7_9_sram;
wire [0:2] sb_mux_size7_9_sram_inv;
wire [0:3] sb_mux_size8_0_sram;
wire [0:3] sb_mux_size8_0_sram_inv;
wire [0:3] sb_mux_size8_10_sram;
wire [0:3] sb_mux_size8_10_sram_inv;
wire [0:3] sb_mux_size8_11_sram;
wire [0:3] sb_mux_size8_11_sram_inv;
wire [0:3] sb_mux_size8_12_sram;
wire [0:3] sb_mux_size8_12_sram_inv;
wire [0:3] sb_mux_size8_13_sram;
wire [0:3] sb_mux_size8_13_sram_inv;
wire [0:3] sb_mux_size8_14_sram;
wire [0:3] sb_mux_size8_14_sram_inv;
wire [0:3] sb_mux_size8_15_sram;
wire [0:3] sb_mux_size8_15_sram_inv;
wire [0:3] sb_mux_size8_1_sram;
wire [0:3] sb_mux_size8_1_sram_inv;
wire [0:3] sb_mux_size8_2_sram;
wire [0:3] sb_mux_size8_2_sram_inv;
wire [0:3] sb_mux_size8_3_sram;
wire [0:3] sb_mux_size8_3_sram_inv;
wire [0:3] sb_mux_size8_4_sram;
wire [0:3] sb_mux_size8_4_sram_inv;
wire [0:3] sb_mux_size8_5_sram;
wire [0:3] sb_mux_size8_5_sram_inv;
wire [0:3] sb_mux_size8_6_sram;
wire [0:3] sb_mux_size8_6_sram_inv;
wire [0:3] sb_mux_size8_7_sram;
wire [0:3] sb_mux_size8_7_sram_inv;
wire [0:3] sb_mux_size8_8_sram;
wire [0:3] sb_mux_size8_8_sram_inv;
wire [0:3] sb_mux_size8_9_sram;
wire [0:3] sb_mux_size8_9_sram_inv;
wire [0:3] sb_mux_size9_0_sram;
wire [0:3] sb_mux_size9_0_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[32] = chanx_right_in[0];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[1];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[2];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[3];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[36] = chanx_right_in[4];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[5];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[6];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[7];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[40] = chanx_right_in[8];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[9];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[10];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[11];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[44] = chanx_right_in[12];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[13];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[14];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[15];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[16];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[17];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[18];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[19];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[52] = chanx_right_in[20];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[21];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[22];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[23];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[56] = chanx_right_in[24];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[25];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[26];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[27];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[60] = chanx_right_in[28];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[29];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[30];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[31];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[0] = chanx_left_in[32];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[33];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[34];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[35];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[4] = chanx_left_in[36];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[37];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[38];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[39];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[8] = chanx_left_in[40];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[41];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[42];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[43];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[12] = chanx_left_in[44];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[45];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[46];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[47];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[16] = chanx_left_in[48];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[49];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[50];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[51];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[20] = chanx_left_in[52];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[53];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[54];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[55];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[24] = chanx_left_in[56];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[57];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[58];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[59];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[28] = chanx_left_in[60];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[61];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[62];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[63];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_[0];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size8 mux_top_track_0 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[0], chanx_left_in[0], chanx_left_in[14], chanx_left_in[28]}),
		.sram(sb_mux_size8_0_sram[0:3]),
		.sram_inv(sb_mux_size8_0_sram_inv[0:3]),
		.out(chany_top_out[0]));

	sb_mux_size8 mux_top_track_24 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chany_bottom_in[15], chanx_left_in[5], chanx_left_in[19]}),
		.sram(sb_mux_size8_1_sram[0:3]),
		.sram_inv(sb_mux_size8_1_sram_inv[0:3]),
		.out(chany_top_out[12]));

	sb_mux_size8 mux_top_track_32 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chany_bottom_in[19], chanx_left_in[4], chanx_left_in[18]}),
		.sram(sb_mux_size8_2_sram[0:3]),
		.sram_inv(sb_mux_size8_2_sram_inv[0:3]),
		.out(chany_top_out[16]));

	sb_mux_size8 mux_top_track_48 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chany_bottom_in[27], chanx_left_in[2], chanx_left_in[16], chanx_left_in[30]}),
		.sram(sb_mux_size8_3_sram[0:3]),
		.sram_inv(sb_mux_size8_3_sram_inv[0:3]),
		.out(chany_top_out[24]));

	sb_mux_size8 mux_top_track_56 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[31], chanx_left_in[1], chanx_left_in[15], chanx_left_in[29]}),
		.sram(sb_mux_size8_4_sram[0:3]),
		.sram_inv(sb_mux_size8_4_sram_inv[0:3]),
		.out(chany_top_out[28]));

	sb_mux_size8 mux_bottom_track_1 (
		.in({chany_top_in[0], bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_left_in[1], chanx_left_in[15], chanx_left_in[29]}),
		.sram(sb_mux_size8_5_sram[0:3]),
		.sram_inv(sb_mux_size8_5_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	sb_mux_size8 mux_bottom_track_3 (
		.in({chany_top_in[1], bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[2], chanx_left_in[16], chanx_left_in[30]}),
		.sram(sb_mux_size8_6_sram[0:3]),
		.sram_inv(sb_mux_size8_6_sram_inv[0:3]),
		.out(chany_bottom_out[1]));

	sb_mux_size8 mux_bottom_track_5 (
		.in({chany_top_in[2], bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chanx_left_in[3], chanx_left_in[17], chanx_left_in[31]}),
		.sram(sb_mux_size8_7_sram[0:3]),
		.sram_inv(sb_mux_size8_7_sram_inv[0:3]),
		.out(chany_bottom_out[2]));

	sb_mux_size8 mux_bottom_track_25 (
		.in({chany_top_in[15], bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chanx_left_in[10], chanx_left_in[24]}),
		.sram(sb_mux_size8_8_sram[0:3]),
		.sram_inv(sb_mux_size8_8_sram_inv[0:3]),
		.out(chany_bottom_out[12]));

	sb_mux_size8 mux_bottom_track_33 (
		.in({chany_top_in[19], bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chanx_left_in[11], chanx_left_in[25]}),
		.sram(sb_mux_size8_9_sram[0:3]),
		.sram_inv(sb_mux_size8_9_sram_inv[0:3]),
		.out(chany_bottom_out[16]));

	sb_mux_size8 mux_bottom_track_41 (
		.in({chany_top_in[23], bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chanx_left_in[12], chanx_left_in[26]}),
		.sram(sb_mux_size8_10_sram[0:3]),
		.sram_inv(sb_mux_size8_10_sram_inv[0:3]),
		.out(chany_bottom_out[20]));

	sb_mux_size8 mux_bottom_track_57 (
		.in({chany_top_in[31], bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chanx_left_in[0], chanx_left_in[14], chanx_left_in[28]}),
		.sram(sb_mux_size8_11_sram[0:3]),
		.sram_inv(sb_mux_size8_11_sram_inv[0:3]),
		.out(chany_bottom_out[28]));

	sb_mux_size8 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[6], chany_bottom_in[6], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_}),
		.sram(sb_mux_size8_12_sram[0:3]),
		.sram_inv(sb_mux_size8_12_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	sb_mux_size8 mux_left_track_3 (
		.in({chany_top_in[8], chany_bottom_in[0], chany_bottom_in[8], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_}),
		.sram(sb_mux_size8_13_sram[0:3]),
		.sram_inv(sb_mux_size8_13_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	sb_mux_size8 mux_left_track_13 (
		.in({chany_top_in[16], chany_bottom_in[5], chany_bottom_in[16], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_}),
		.sram(sb_mux_size8_14_sram[0:3]),
		.sram_inv(sb_mux_size8_14_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	sb_mux_size8 mux_left_track_15 (
		.in({chany_top_in[17], chany_bottom_in[7], chany_bottom_in[17], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_}),
		.sram(sb_mux_size8_15_sram[0:3]),
		.sram_inv(sb_mux_size8_15_sram_inv[0:3]),
		.out(chanx_left_out[7]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_0 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[0:3]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[0:3]),
		.mem_out(sb_mux_size8_0_sram[0:3]),
		.mem_outb(sb_mux_size8_0_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_24 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[31:34]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[31:34]),
		.mem_out(sb_mux_size8_1_sram[0:3]),
		.mem_outb(sb_mux_size8_1_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_32 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[35:38]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[35:38]),
		.mem_out(sb_mux_size8_2_sram[0:3]),
		.mem_outb(sb_mux_size8_2_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_48 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[43:46]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[43:46]),
		.mem_out(sb_mux_size8_3_sram[0:3]),
		.mem_outb(sb_mux_size8_3_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_top_track_56 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[47:50]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[47:50]),
		.mem_out(sb_mux_size8_4_sram[0:3]),
		.mem_outb(sb_mux_size8_4_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_1 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[115:118]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[115:118]),
		.mem_out(sb_mux_size8_5_sram[0:3]),
		.mem_outb(sb_mux_size8_5_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_3 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[119:122]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[119:122]),
		.mem_out(sb_mux_size8_6_sram[0:3]),
		.mem_outb(sb_mux_size8_6_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_5 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[123:126]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[123:126]),
		.mem_out(sb_mux_size8_7_sram[0:3]),
		.mem_outb(sb_mux_size8_7_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_25 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[148:151]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[148:151]),
		.mem_out(sb_mux_size8_8_sram[0:3]),
		.mem_outb(sb_mux_size8_8_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_33 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[152:155]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[152:155]),
		.mem_out(sb_mux_size8_9_sram[0:3]),
		.mem_outb(sb_mux_size8_9_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_41 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[156:159]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[156:159]),
		.mem_out(sb_mux_size8_10_sram[0:3]),
		.mem_outb(sb_mux_size8_10_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_bottom_track_57 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[163:166]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[163:166]),
		.mem_out(sb_mux_size8_11_sram[0:3]),
		.mem_outb(sb_mux_size8_11_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_1 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[231:234]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[231:234]),
		.mem_out(sb_mux_size8_12_sram[0:3]),
		.mem_outb(sb_mux_size8_12_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_3 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[235:238]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[235:238]),
		.mem_out(sb_mux_size8_13_sram[0:3]),
		.mem_outb(sb_mux_size8_13_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_13 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[251:254]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[251:254]),
		.mem_out(sb_mux_size8_14_sram[0:3]),
		.mem_outb(sb_mux_size8_14_sram_inv[0:3]));

	sb_mux_size8_feedthrough_mem feedthrough_mem_left_track_15 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[255:258]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[255:258]),
		.mem_out(sb_mux_size8_15_sram[0:3]),
		.mem_outb(sb_mux_size8_15_sram_inv[0:3]));

	sb_mux_size7 mux_top_track_2 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, chany_bottom_in[1], chanx_left_in[13], chanx_left_in[27]}),
		.sram(sb_mux_size7_0_sram[0:2]),
		.sram_inv(sb_mux_size7_0_sram_inv[0:2]),
		.out(chany_top_out[1]));

	sb_mux_size7 mux_top_track_4 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chany_bottom_in[2], chanx_left_in[12], chanx_left_in[26]}),
		.sram(sb_mux_size7_1_sram[0:2]),
		.sram_inv(sb_mux_size7_1_sram_inv[0:2]),
		.out(chany_top_out[2]));

	sb_mux_size7 mux_top_track_6 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chany_bottom_in[3], chanx_left_in[11], chanx_left_in[25]}),
		.sram(sb_mux_size7_2_sram[0:2]),
		.sram_inv(sb_mux_size7_2_sram_inv[0:2]),
		.out(chany_top_out[3]));

	sb_mux_size7 mux_top_track_8 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chany_bottom_in[4], chanx_left_in[10], chanx_left_in[24]}),
		.sram(sb_mux_size7_3_sram[0:2]),
		.sram_inv(sb_mux_size7_3_sram_inv[0:2]),
		.out(chany_top_out[4]));

	sb_mux_size7 mux_bottom_track_7 (
		.in({chany_top_in[3], bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chanx_left_in[4], chanx_left_in[18]}),
		.sram(sb_mux_size7_4_sram[0:2]),
		.sram_inv(sb_mux_size7_4_sram_inv[0:2]),
		.out(chany_bottom_out[3]));

	sb_mux_size7 mux_bottom_track_9 (
		.in({chany_top_in[4], bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chanx_left_in[5], chanx_left_in[19]}),
		.sram(sb_mux_size7_5_sram[0:2]),
		.sram_inv(sb_mux_size7_5_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	sb_mux_size7 mux_bottom_track_49 (
		.in({chany_top_in[27], bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, chanx_left_in[13], chanx_left_in[27]}),
		.sram(sb_mux_size7_6_sram[0:2]),
		.sram_inv(sb_mux_size7_6_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	sb_mux_size7 mux_left_track_5 (
		.in({chany_top_in[10], chany_bottom_in[1], chany_bottom_in[10], left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_}),
		.sram(sb_mux_size7_7_sram[0:2]),
		.sram_inv(sb_mux_size7_7_sram_inv[0:2]),
		.out(chanx_left_out[2]));

	sb_mux_size7 mux_left_track_7 (
		.in({chany_top_in[12], chany_bottom_in[2], chany_bottom_in[12], left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_}),
		.sram(sb_mux_size7_8_sram[0:2]),
		.sram_inv(sb_mux_size7_8_sram_inv[0:2]),
		.out(chanx_left_out[3]));

	sb_mux_size7 mux_left_track_9 (
		.in({chany_top_in[13], chany_bottom_in[3], chany_bottom_in[13], left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_}),
		.sram(sb_mux_size7_9_sram[0:2]),
		.sram_inv(sb_mux_size7_9_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	sb_mux_size7 mux_left_track_11 (
		.in({chany_top_in[14], chany_bottom_in[4], chany_bottom_in[14], left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_}),
		.sram(sb_mux_size7_10_sram[0:2]),
		.sram_inv(sb_mux_size7_10_sram_inv[0:2]),
		.out(chanx_left_out[5]));

	sb_mux_size7 mux_left_track_17 (
		.in({chany_top_in[18], chany_bottom_in[9], chany_bottom_in[18], left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_}),
		.sram(sb_mux_size7_11_sram[0:2]),
		.sram_inv(sb_mux_size7_11_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	sb_mux_size7 mux_left_track_19 (
		.in({chany_top_in[20], chany_bottom_in[11], chany_bottom_in[20], left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_}),
		.sram(sb_mux_size7_12_sram[0:2]),
		.sram_inv(sb_mux_size7_12_sram_inv[0:2]),
		.out(chanx_left_out[9]));

	sb_mux_size7 mux_left_track_21 (
		.in({chany_top_in[21], chany_bottom_in[15], chany_bottom_in[21], left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_}),
		.sram(sb_mux_size7_13_sram[0:2]),
		.sram_inv(sb_mux_size7_13_sram_inv[0:2]),
		.out(chanx_left_out[10]));

	sb_mux_size7 mux_left_track_23 (
		.in({chany_top_in[22], chany_bottom_in[19], chany_bottom_in[22], left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_}),
		.sram(sb_mux_size7_14_sram[0:2]),
		.sram_inv(sb_mux_size7_14_sram_inv[0:2]),
		.out(chanx_left_out[11]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_2 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[4:6]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[4:6]),
		.mem_out(sb_mux_size7_0_sram[0:2]),
		.mem_outb(sb_mux_size7_0_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_4 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[7:9]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[7:9]),
		.mem_out(sb_mux_size7_1_sram[0:2]),
		.mem_outb(sb_mux_size7_1_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_6 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[10:12]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[10:12]),
		.mem_out(sb_mux_size7_2_sram[0:2]),
		.mem_outb(sb_mux_size7_2_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_top_track_8 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[13:15]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[13:15]),
		.mem_out(sb_mux_size7_3_sram[0:2]),
		.mem_outb(sb_mux_size7_3_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_7 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[127:129]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[127:129]),
		.mem_out(sb_mux_size7_4_sram[0:2]),
		.mem_outb(sb_mux_size7_4_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_9 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[130:132]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[130:132]),
		.mem_out(sb_mux_size7_5_sram[0:2]),
		.mem_outb(sb_mux_size7_5_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_bottom_track_49 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[160:162]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[160:162]),
		.mem_out(sb_mux_size7_6_sram[0:2]),
		.mem_outb(sb_mux_size7_6_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_5 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[239:241]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[239:241]),
		.mem_out(sb_mux_size7_7_sram[0:2]),
		.mem_outb(sb_mux_size7_7_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_7 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[242:244]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[242:244]),
		.mem_out(sb_mux_size7_8_sram[0:2]),
		.mem_outb(sb_mux_size7_8_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_9 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[245:247]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[245:247]),
		.mem_out(sb_mux_size7_9_sram[0:2]),
		.mem_outb(sb_mux_size7_9_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_11 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[248:250]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[248:250]),
		.mem_out(sb_mux_size7_10_sram[0:2]),
		.mem_outb(sb_mux_size7_10_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_17 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[259:261]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[259:261]),
		.mem_out(sb_mux_size7_11_sram[0:2]),
		.mem_outb(sb_mux_size7_11_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_19 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[262:264]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[262:264]),
		.mem_out(sb_mux_size7_12_sram[0:2]),
		.mem_outb(sb_mux_size7_12_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_21 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[265:267]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[265:267]),
		.mem_out(sb_mux_size7_13_sram[0:2]),
		.mem_outb(sb_mux_size7_13_sram_inv[0:2]));

	sb_mux_size7_feedthrough_mem feedthrough_mem_left_track_23 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[268:270]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[268:270]),
		.mem_out(sb_mux_size7_14_sram[0:2]),
		.mem_outb(sb_mux_size7_14_sram_inv[0:2]));

	sb_mux_size6 mux_top_track_10 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chany_bottom_in[5], chanx_left_in[9], chanx_left_in[23]}),
		.sram(sb_mux_size6_0_sram[0:2]),
		.sram_inv(sb_mux_size6_0_sram_inv[0:2]),
		.out(chany_top_out[5]));

	sb_mux_size6 mux_bottom_track_11 (
		.in({chany_top_in[5], bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, chanx_left_in[6], chanx_left_in[20]}),
		.sram(sb_mux_size6_1_sram[0:2]),
		.sram_inv(sb_mux_size6_1_sram_inv[0:2]),
		.out(chany_bottom_out[5]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_top_track_10 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[16:18]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[16:18]),
		.mem_out(sb_mux_size6_0_sram[0:2]),
		.mem_outb(sb_mux_size6_0_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_bottom_track_11 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[133:135]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[133:135]),
		.mem_out(sb_mux_size6_1_sram[0:2]),
		.mem_outb(sb_mux_size6_1_sram_inv[0:2]));

	sb_mux_size11 mux_top_track_12 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chany_bottom_in[7], chanx_left_in[8], chanx_left_in[22]}),
		.sram(sb_mux_size11_0_sram[0:3]),
		.sram_inv(sb_mux_size11_0_sram_inv[0:3]),
		.out(chany_top_out[6]));

	sb_mux_size11 mux_top_track_16 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chany_bottom_in[9], chanx_left_in[7], chanx_left_in[21]}),
		.sram(sb_mux_size11_1_sram[0:3]),
		.sram_inv(sb_mux_size11_1_sram_inv[0:3]),
		.out(chany_top_out[8]));

	sb_mux_size11 mux_bottom_track_13 (
		.in({chany_top_in[7], bottom_right_grid_left_width_0_height_0_subtile_0__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_match0_o_0_, chanx_left_in[7], chanx_left_in[21]}),
		.sram(sb_mux_size11_2_sram[0:3]),
		.sram_inv(sb_mux_size11_2_sram_inv[0:3]),
		.out(chany_bottom_out[6]));

	sb_mux_size11 mux_bottom_track_17 (
		.in({chany_top_in[9], bottom_right_grid_left_width_0_height_0_subtile_1__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_2_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chanx_left_in[8], chanx_left_in[22]}),
		.sram(sb_mux_size11_3_sram[0:3]),
		.sram_inv(sb_mux_size11_3_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_top_track_12 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[19:22]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[19:22]),
		.mem_out(sb_mux_size11_0_sram[0:3]),
		.mem_outb(sb_mux_size11_0_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_top_track_16 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[23:26]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[23:26]),
		.mem_out(sb_mux_size11_1_sram[0:3]),
		.mem_outb(sb_mux_size11_1_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_bottom_track_13 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[136:139]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[136:139]),
		.mem_out(sb_mux_size11_2_sram[0:3]),
		.mem_outb(sb_mux_size11_2_sram_inv[0:3]));

	sb_mux_size11_feedthrough_mem feedthrough_mem_bottom_track_17 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[140:143]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[140:143]),
		.mem_out(sb_mux_size11_3_sram[0:3]),
		.mem_outb(sb_mux_size11_3_sram_inv[0:3]));

	sb_mux_size10 mux_top_track_20 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chany_bottom_in[11], chanx_left_in[6], chanx_left_in[20]}),
		.sram(sb_mux_size10_0_sram[0:3]),
		.sram_inv(sb_mux_size10_0_sram_inv[0:3]),
		.out(chany_top_out[10]));

	sb_mux_size10 mux_bottom_track_21 (
		.in({chany_top_in[11], bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_6_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_match0_o_0_, chanx_left_in[9], chanx_left_in[23]}),
		.sram(sb_mux_size10_1_sram[0:3]),
		.sram_inv(sb_mux_size10_1_sram_inv[0:3]),
		.out(chany_bottom_out[10]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_top_track_20 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[27:30]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[27:30]),
		.mem_out(sb_mux_size10_0_sram[0:3]),
		.mem_outb(sb_mux_size10_0_sram_inv[0:3]));

	sb_mux_size10_feedthrough_mem feedthrough_mem_bottom_track_21 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[144:147]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[144:147]),
		.mem_out(sb_mux_size10_1_sram[0:3]),
		.mem_outb(sb_mux_size10_1_sram_inv[0:3]));

	sb_mux_size9 mux_top_track_40 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_a2f_o_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_a2f_o_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_4_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_match0_o_0_, chany_bottom_in[23], chanx_left_in[3], chanx_left_in[17], chanx_left_in[31]}),
		.sram(sb_mux_size9_0_sram[0:3]),
		.sram_inv(sb_mux_size9_0_sram_inv[0:3]),
		.out(chany_top_out[20]));

	sb_mux_size9_feedthrough_mem feedthrough_mem_top_track_40 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[39:42]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[39:42]),
		.mem_out(sb_mux_size9_0_sram[0:3]),
		.mem_outb(sb_mux_size9_0_sram_inv[0:3]));

	clk_mux_size3 mux_top_track_64 (
		.in({chanx_right_in[0], chany_bottom_in[32], chanx_left_in[32]}),
		.sram(clk_mux_size3_0_sram[0:1]),
		.sram_inv(clk_mux_size3_0_sram_inv[0:1]),
		.out(chany_top_out[32]));

	clk_mux_size3 mux_top_track_66 (
		.in({chanx_right_in[1], chany_bottom_in[33], chanx_left_in[33]}),
		.sram(clk_mux_size3_1_sram[0:1]),
		.sram_inv(clk_mux_size3_1_sram_inv[0:1]),
		.out(chany_top_out[33]));

	clk_mux_size3 mux_top_track_68 (
		.in({chanx_right_in[2], chany_bottom_in[34], chanx_left_in[34]}),
		.sram(clk_mux_size3_2_sram[0:1]),
		.sram_inv(clk_mux_size3_2_sram_inv[0:1]),
		.out(chany_top_out[34]));

	clk_mux_size3 mux_top_track_70 (
		.in({chanx_right_in[3], chany_bottom_in[35], chanx_left_in[35]}),
		.sram(clk_mux_size3_3_sram[0:1]),
		.sram_inv(clk_mux_size3_3_sram_inv[0:1]),
		.out(chany_top_out[35]));

	clk_mux_size3 mux_top_track_72 (
		.in({chanx_right_in[4], chany_bottom_in[36], chanx_left_in[36]}),
		.sram(clk_mux_size3_4_sram[0:1]),
		.sram_inv(clk_mux_size3_4_sram_inv[0:1]),
		.out(chany_top_out[36]));

	clk_mux_size3 mux_top_track_74 (
		.in({chanx_right_in[5], chany_bottom_in[37], chanx_left_in[37]}),
		.sram(clk_mux_size3_5_sram[0:1]),
		.sram_inv(clk_mux_size3_5_sram_inv[0:1]),
		.out(chany_top_out[37]));

	clk_mux_size3 mux_top_track_76 (
		.in({chanx_right_in[6], chany_bottom_in[38], chanx_left_in[38]}),
		.sram(clk_mux_size3_6_sram[0:1]),
		.sram_inv(clk_mux_size3_6_sram_inv[0:1]),
		.out(chany_top_out[38]));

	clk_mux_size3 mux_top_track_78 (
		.in({chanx_right_in[7], chany_bottom_in[39], chanx_left_in[39]}),
		.sram(clk_mux_size3_7_sram[0:1]),
		.sram_inv(clk_mux_size3_7_sram_inv[0:1]),
		.out(chany_top_out[39]));

	clk_mux_size3 mux_top_track_80 (
		.in({chanx_right_in[8], chany_bottom_in[40], chanx_left_in[40]}),
		.sram(clk_mux_size3_8_sram[0:1]),
		.sram_inv(clk_mux_size3_8_sram_inv[0:1]),
		.out(chany_top_out[40]));

	clk_mux_size3 mux_top_track_82 (
		.in({chanx_right_in[9], chany_bottom_in[41], chanx_left_in[41]}),
		.sram(clk_mux_size3_9_sram[0:1]),
		.sram_inv(clk_mux_size3_9_sram_inv[0:1]),
		.out(chany_top_out[41]));

	clk_mux_size3 mux_top_track_84 (
		.in({chanx_right_in[10], chany_bottom_in[42], chanx_left_in[42]}),
		.sram(clk_mux_size3_10_sram[0:1]),
		.sram_inv(clk_mux_size3_10_sram_inv[0:1]),
		.out(chany_top_out[42]));

	clk_mux_size3 mux_top_track_86 (
		.in({chanx_right_in[11], chany_bottom_in[43], chanx_left_in[43]}),
		.sram(clk_mux_size3_11_sram[0:1]),
		.sram_inv(clk_mux_size3_11_sram_inv[0:1]),
		.out(chany_top_out[43]));

	clk_mux_size3 mux_top_track_88 (
		.in({chanx_right_in[12], chany_bottom_in[44], chanx_left_in[44]}),
		.sram(clk_mux_size3_12_sram[0:1]),
		.sram_inv(clk_mux_size3_12_sram_inv[0:1]),
		.out(chany_top_out[44]));

	clk_mux_size3 mux_top_track_90 (
		.in({chanx_right_in[13], chany_bottom_in[45], chanx_left_in[45]}),
		.sram(clk_mux_size3_13_sram[0:1]),
		.sram_inv(clk_mux_size3_13_sram_inv[0:1]),
		.out(chany_top_out[45]));

	clk_mux_size3 mux_top_track_92 (
		.in({chanx_right_in[14], chany_bottom_in[46], chanx_left_in[46]}),
		.sram(clk_mux_size3_14_sram[0:1]),
		.sram_inv(clk_mux_size3_14_sram_inv[0:1]),
		.out(chany_top_out[46]));

	clk_mux_size3 mux_top_track_94 (
		.in({chanx_right_in[15], chany_bottom_in[47], chanx_left_in[47]}),
		.sram(clk_mux_size3_15_sram[0:1]),
		.sram_inv(clk_mux_size3_15_sram_inv[0:1]),
		.out(chany_top_out[47]));

	clk_mux_size3 mux_top_track_96 (
		.in({chanx_right_in[16], chany_bottom_in[48], chanx_left_in[48]}),
		.sram(clk_mux_size3_16_sram[0:1]),
		.sram_inv(clk_mux_size3_16_sram_inv[0:1]),
		.out(chany_top_out[48]));

	clk_mux_size3 mux_top_track_98 (
		.in({chanx_right_in[17], chany_bottom_in[49], chanx_left_in[49]}),
		.sram(clk_mux_size3_17_sram[0:1]),
		.sram_inv(clk_mux_size3_17_sram_inv[0:1]),
		.out(chany_top_out[49]));

	clk_mux_size3 mux_top_track_100 (
		.in({chanx_right_in[18], chany_bottom_in[50], chanx_left_in[50]}),
		.sram(clk_mux_size3_18_sram[0:1]),
		.sram_inv(clk_mux_size3_18_sram_inv[0:1]),
		.out(chany_top_out[50]));

	clk_mux_size3 mux_top_track_102 (
		.in({chanx_right_in[19], chany_bottom_in[51], chanx_left_in[51]}),
		.sram(clk_mux_size3_19_sram[0:1]),
		.sram_inv(clk_mux_size3_19_sram_inv[0:1]),
		.out(chany_top_out[51]));

	clk_mux_size3 mux_top_track_104 (
		.in({chanx_right_in[20], chany_bottom_in[52], chanx_left_in[52]}),
		.sram(clk_mux_size3_20_sram[0:1]),
		.sram_inv(clk_mux_size3_20_sram_inv[0:1]),
		.out(chany_top_out[52]));

	clk_mux_size3 mux_top_track_106 (
		.in({chanx_right_in[21], chany_bottom_in[53], chanx_left_in[53]}),
		.sram(clk_mux_size3_21_sram[0:1]),
		.sram_inv(clk_mux_size3_21_sram_inv[0:1]),
		.out(chany_top_out[53]));

	clk_mux_size3 mux_top_track_108 (
		.in({chanx_right_in[22], chany_bottom_in[54], chanx_left_in[54]}),
		.sram(clk_mux_size3_22_sram[0:1]),
		.sram_inv(clk_mux_size3_22_sram_inv[0:1]),
		.out(chany_top_out[54]));

	clk_mux_size3 mux_top_track_110 (
		.in({chanx_right_in[23], chany_bottom_in[55], chanx_left_in[55]}),
		.sram(clk_mux_size3_23_sram[0:1]),
		.sram_inv(clk_mux_size3_23_sram_inv[0:1]),
		.out(chany_top_out[55]));

	clk_mux_size3 mux_top_track_112 (
		.in({chanx_right_in[24], chany_bottom_in[56], chanx_left_in[56]}),
		.sram(clk_mux_size3_24_sram[0:1]),
		.sram_inv(clk_mux_size3_24_sram_inv[0:1]),
		.out(chany_top_out[56]));

	clk_mux_size3 mux_top_track_114 (
		.in({chanx_right_in[25], chany_bottom_in[57], chanx_left_in[57]}),
		.sram(clk_mux_size3_25_sram[0:1]),
		.sram_inv(clk_mux_size3_25_sram_inv[0:1]),
		.out(chany_top_out[57]));

	clk_mux_size3 mux_top_track_116 (
		.in({chanx_right_in[26], chany_bottom_in[58], chanx_left_in[58]}),
		.sram(clk_mux_size3_26_sram[0:1]),
		.sram_inv(clk_mux_size3_26_sram_inv[0:1]),
		.out(chany_top_out[58]));

	clk_mux_size3 mux_top_track_118 (
		.in({chanx_right_in[27], chany_bottom_in[59], chanx_left_in[59]}),
		.sram(clk_mux_size3_27_sram[0:1]),
		.sram_inv(clk_mux_size3_27_sram_inv[0:1]),
		.out(chany_top_out[59]));

	clk_mux_size3 mux_top_track_120 (
		.in({chanx_right_in[28], chany_bottom_in[60], chanx_left_in[60]}),
		.sram(clk_mux_size3_28_sram[0:1]),
		.sram_inv(clk_mux_size3_28_sram_inv[0:1]),
		.out(chany_top_out[60]));

	clk_mux_size3 mux_top_track_122 (
		.in({chanx_right_in[29], chany_bottom_in[61], chanx_left_in[61]}),
		.sram(clk_mux_size3_29_sram[0:1]),
		.sram_inv(clk_mux_size3_29_sram_inv[0:1]),
		.out(chany_top_out[61]));

	clk_mux_size3 mux_top_track_124 (
		.in({chanx_right_in[30], chany_bottom_in[62], chanx_left_in[62]}),
		.sram(clk_mux_size3_30_sram[0:1]),
		.sram_inv(clk_mux_size3_30_sram_inv[0:1]),
		.out(chany_top_out[62]));

	clk_mux_size3 mux_top_track_126 (
		.in({chanx_right_in[31], chany_bottom_in[63], chanx_left_in[63]}),
		.sram(clk_mux_size3_31_sram[0:1]),
		.sram_inv(clk_mux_size3_31_sram_inv[0:1]),
		.out(chany_top_out[63]));

	clk_mux_size3 mux_bottom_track_65 (
		.in({chany_top_in[32], chanx_right_in[0], chanx_left_in[32]}),
		.sram(clk_mux_size3_32_sram[0:1]),
		.sram_inv(clk_mux_size3_32_sram_inv[0:1]),
		.out(chany_bottom_out[32]));

	clk_mux_size3 mux_bottom_track_67 (
		.in({chany_top_in[33], chanx_right_in[1], chanx_left_in[33]}),
		.sram(clk_mux_size3_33_sram[0:1]),
		.sram_inv(clk_mux_size3_33_sram_inv[0:1]),
		.out(chany_bottom_out[33]));

	clk_mux_size3 mux_bottom_track_69 (
		.in({chany_top_in[34], chanx_right_in[2], chanx_left_in[34]}),
		.sram(clk_mux_size3_34_sram[0:1]),
		.sram_inv(clk_mux_size3_34_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	clk_mux_size3 mux_bottom_track_71 (
		.in({chany_top_in[35], chanx_right_in[3], chanx_left_in[35]}),
		.sram(clk_mux_size3_35_sram[0:1]),
		.sram_inv(clk_mux_size3_35_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	clk_mux_size3 mux_bottom_track_73 (
		.in({chany_top_in[36], chanx_right_in[4], chanx_left_in[36]}),
		.sram(clk_mux_size3_36_sram[0:1]),
		.sram_inv(clk_mux_size3_36_sram_inv[0:1]),
		.out(chany_bottom_out[36]));

	clk_mux_size3 mux_bottom_track_75 (
		.in({chany_top_in[37], chanx_right_in[5], chanx_left_in[37]}),
		.sram(clk_mux_size3_37_sram[0:1]),
		.sram_inv(clk_mux_size3_37_sram_inv[0:1]),
		.out(chany_bottom_out[37]));

	clk_mux_size3 mux_bottom_track_77 (
		.in({chany_top_in[38], chanx_right_in[6], chanx_left_in[38]}),
		.sram(clk_mux_size3_38_sram[0:1]),
		.sram_inv(clk_mux_size3_38_sram_inv[0:1]),
		.out(chany_bottom_out[38]));

	clk_mux_size3 mux_bottom_track_79 (
		.in({chany_top_in[39], chanx_right_in[7], chanx_left_in[39]}),
		.sram(clk_mux_size3_39_sram[0:1]),
		.sram_inv(clk_mux_size3_39_sram_inv[0:1]),
		.out(chany_bottom_out[39]));

	clk_mux_size3 mux_bottom_track_81 (
		.in({chany_top_in[40], chanx_right_in[8], chanx_left_in[40]}),
		.sram(clk_mux_size3_40_sram[0:1]),
		.sram_inv(clk_mux_size3_40_sram_inv[0:1]),
		.out(chany_bottom_out[40]));

	clk_mux_size3 mux_bottom_track_83 (
		.in({chany_top_in[41], chanx_right_in[9], chanx_left_in[41]}),
		.sram(clk_mux_size3_41_sram[0:1]),
		.sram_inv(clk_mux_size3_41_sram_inv[0:1]),
		.out(chany_bottom_out[41]));

	clk_mux_size3 mux_bottom_track_85 (
		.in({chany_top_in[42], chanx_right_in[10], chanx_left_in[42]}),
		.sram(clk_mux_size3_42_sram[0:1]),
		.sram_inv(clk_mux_size3_42_sram_inv[0:1]),
		.out(chany_bottom_out[42]));

	clk_mux_size3 mux_bottom_track_87 (
		.in({chany_top_in[43], chanx_right_in[11], chanx_left_in[43]}),
		.sram(clk_mux_size3_43_sram[0:1]),
		.sram_inv(clk_mux_size3_43_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	clk_mux_size3 mux_bottom_track_89 (
		.in({chany_top_in[44], chanx_right_in[12], chanx_left_in[44]}),
		.sram(clk_mux_size3_44_sram[0:1]),
		.sram_inv(clk_mux_size3_44_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	clk_mux_size3 mux_bottom_track_91 (
		.in({chany_top_in[45], chanx_right_in[13], chanx_left_in[45]}),
		.sram(clk_mux_size3_45_sram[0:1]),
		.sram_inv(clk_mux_size3_45_sram_inv[0:1]),
		.out(chany_bottom_out[45]));

	clk_mux_size3 mux_bottom_track_93 (
		.in({chany_top_in[46], chanx_right_in[14], chanx_left_in[46]}),
		.sram(clk_mux_size3_46_sram[0:1]),
		.sram_inv(clk_mux_size3_46_sram_inv[0:1]),
		.out(chany_bottom_out[46]));

	clk_mux_size3 mux_bottom_track_95 (
		.in({chany_top_in[47], chanx_right_in[15], chanx_left_in[47]}),
		.sram(clk_mux_size3_47_sram[0:1]),
		.sram_inv(clk_mux_size3_47_sram_inv[0:1]),
		.out(chany_bottom_out[47]));

	clk_mux_size3 mux_bottom_track_97 (
		.in({chany_top_in[48], chanx_right_in[16], chanx_left_in[48]}),
		.sram(clk_mux_size3_48_sram[0:1]),
		.sram_inv(clk_mux_size3_48_sram_inv[0:1]),
		.out(chany_bottom_out[48]));

	clk_mux_size3 mux_bottom_track_99 (
		.in({chany_top_in[49], chanx_right_in[17], chanx_left_in[49]}),
		.sram(clk_mux_size3_49_sram[0:1]),
		.sram_inv(clk_mux_size3_49_sram_inv[0:1]),
		.out(chany_bottom_out[49]));

	clk_mux_size3 mux_bottom_track_101 (
		.in({chany_top_in[50], chanx_right_in[18], chanx_left_in[50]}),
		.sram(clk_mux_size3_50_sram[0:1]),
		.sram_inv(clk_mux_size3_50_sram_inv[0:1]),
		.out(chany_bottom_out[50]));

	clk_mux_size3 mux_bottom_track_103 (
		.in({chany_top_in[51], chanx_right_in[19], chanx_left_in[51]}),
		.sram(clk_mux_size3_51_sram[0:1]),
		.sram_inv(clk_mux_size3_51_sram_inv[0:1]),
		.out(chany_bottom_out[51]));

	clk_mux_size3 mux_bottom_track_105 (
		.in({chany_top_in[52], chanx_right_in[20], chanx_left_in[52]}),
		.sram(clk_mux_size3_52_sram[0:1]),
		.sram_inv(clk_mux_size3_52_sram_inv[0:1]),
		.out(chany_bottom_out[52]));

	clk_mux_size3 mux_bottom_track_107 (
		.in({chany_top_in[53], chanx_right_in[21], chanx_left_in[53]}),
		.sram(clk_mux_size3_53_sram[0:1]),
		.sram_inv(clk_mux_size3_53_sram_inv[0:1]),
		.out(chany_bottom_out[53]));

	clk_mux_size3 mux_bottom_track_109 (
		.in({chany_top_in[54], chanx_right_in[22], chanx_left_in[54]}),
		.sram(clk_mux_size3_54_sram[0:1]),
		.sram_inv(clk_mux_size3_54_sram_inv[0:1]),
		.out(chany_bottom_out[54]));

	clk_mux_size3 mux_bottom_track_111 (
		.in({chany_top_in[55], chanx_right_in[23], chanx_left_in[55]}),
		.sram(clk_mux_size3_55_sram[0:1]),
		.sram_inv(clk_mux_size3_55_sram_inv[0:1]),
		.out(chany_bottom_out[55]));

	clk_mux_size3 mux_bottom_track_113 (
		.in({chany_top_in[56], chanx_right_in[24], chanx_left_in[56]}),
		.sram(clk_mux_size3_56_sram[0:1]),
		.sram_inv(clk_mux_size3_56_sram_inv[0:1]),
		.out(chany_bottom_out[56]));

	clk_mux_size3 mux_bottom_track_115 (
		.in({chany_top_in[57], chanx_right_in[25], chanx_left_in[57]}),
		.sram(clk_mux_size3_57_sram[0:1]),
		.sram_inv(clk_mux_size3_57_sram_inv[0:1]),
		.out(chany_bottom_out[57]));

	clk_mux_size3 mux_bottom_track_117 (
		.in({chany_top_in[58], chanx_right_in[26], chanx_left_in[58]}),
		.sram(clk_mux_size3_58_sram[0:1]),
		.sram_inv(clk_mux_size3_58_sram_inv[0:1]),
		.out(chany_bottom_out[58]));

	clk_mux_size3 mux_bottom_track_119 (
		.in({chany_top_in[59], chanx_right_in[27], chanx_left_in[59]}),
		.sram(clk_mux_size3_59_sram[0:1]),
		.sram_inv(clk_mux_size3_59_sram_inv[0:1]),
		.out(chany_bottom_out[59]));

	clk_mux_size3 mux_bottom_track_121 (
		.in({chany_top_in[60], chanx_right_in[28], chanx_left_in[60]}),
		.sram(clk_mux_size3_60_sram[0:1]),
		.sram_inv(clk_mux_size3_60_sram_inv[0:1]),
		.out(chany_bottom_out[60]));

	clk_mux_size3 mux_bottom_track_123 (
		.in({chany_top_in[61], chanx_right_in[29], chanx_left_in[61]}),
		.sram(clk_mux_size3_61_sram[0:1]),
		.sram_inv(clk_mux_size3_61_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	clk_mux_size3 mux_bottom_track_125 (
		.in({chany_top_in[62], chanx_right_in[30], chanx_left_in[62]}),
		.sram(clk_mux_size3_62_sram[0:1]),
		.sram_inv(clk_mux_size3_62_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	clk_mux_size3 mux_bottom_track_127 (
		.in({chany_top_in[63], chanx_right_in[31], chanx_left_in[63]}),
		.sram(clk_mux_size3_63_sram[0:1]),
		.sram_inv(clk_mux_size3_63_sram_inv[0:1]),
		.out(chany_bottom_out[63]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_64 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[51:52]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[51:52]),
		.mem_out(clk_mux_size3_0_sram[0:1]),
		.mem_outb(clk_mux_size3_0_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_66 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[53:54]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[53:54]),
		.mem_out(clk_mux_size3_1_sram[0:1]),
		.mem_outb(clk_mux_size3_1_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_68 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[55:56]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[55:56]),
		.mem_out(clk_mux_size3_2_sram[0:1]),
		.mem_outb(clk_mux_size3_2_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_70 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[57:58]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[57:58]),
		.mem_out(clk_mux_size3_3_sram[0:1]),
		.mem_outb(clk_mux_size3_3_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_72 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[59:60]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[59:60]),
		.mem_out(clk_mux_size3_4_sram[0:1]),
		.mem_outb(clk_mux_size3_4_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_74 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[61:62]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[61:62]),
		.mem_out(clk_mux_size3_5_sram[0:1]),
		.mem_outb(clk_mux_size3_5_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_76 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[63:64]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[63:64]),
		.mem_out(clk_mux_size3_6_sram[0:1]),
		.mem_outb(clk_mux_size3_6_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_78 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[65:66]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[65:66]),
		.mem_out(clk_mux_size3_7_sram[0:1]),
		.mem_outb(clk_mux_size3_7_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_80 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[67:68]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[67:68]),
		.mem_out(clk_mux_size3_8_sram[0:1]),
		.mem_outb(clk_mux_size3_8_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_82 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[69:70]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[69:70]),
		.mem_out(clk_mux_size3_9_sram[0:1]),
		.mem_outb(clk_mux_size3_9_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_84 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[71:72]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[71:72]),
		.mem_out(clk_mux_size3_10_sram[0:1]),
		.mem_outb(clk_mux_size3_10_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_86 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[73:74]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[73:74]),
		.mem_out(clk_mux_size3_11_sram[0:1]),
		.mem_outb(clk_mux_size3_11_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_88 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[75:76]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[75:76]),
		.mem_out(clk_mux_size3_12_sram[0:1]),
		.mem_outb(clk_mux_size3_12_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_90 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[77:78]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[77:78]),
		.mem_out(clk_mux_size3_13_sram[0:1]),
		.mem_outb(clk_mux_size3_13_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_92 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[79:80]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[79:80]),
		.mem_out(clk_mux_size3_14_sram[0:1]),
		.mem_outb(clk_mux_size3_14_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_94 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[81:82]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[81:82]),
		.mem_out(clk_mux_size3_15_sram[0:1]),
		.mem_outb(clk_mux_size3_15_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_96 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[83:84]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[83:84]),
		.mem_out(clk_mux_size3_16_sram[0:1]),
		.mem_outb(clk_mux_size3_16_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_98 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[85:86]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[85:86]),
		.mem_out(clk_mux_size3_17_sram[0:1]),
		.mem_outb(clk_mux_size3_17_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_100 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[87:88]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[87:88]),
		.mem_out(clk_mux_size3_18_sram[0:1]),
		.mem_outb(clk_mux_size3_18_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_102 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[89:90]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[89:90]),
		.mem_out(clk_mux_size3_19_sram[0:1]),
		.mem_outb(clk_mux_size3_19_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_104 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[91:92]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[91:92]),
		.mem_out(clk_mux_size3_20_sram[0:1]),
		.mem_outb(clk_mux_size3_20_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_106 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[93:94]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[93:94]),
		.mem_out(clk_mux_size3_21_sram[0:1]),
		.mem_outb(clk_mux_size3_21_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_108 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[95:96]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[95:96]),
		.mem_out(clk_mux_size3_22_sram[0:1]),
		.mem_outb(clk_mux_size3_22_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_110 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[97:98]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[97:98]),
		.mem_out(clk_mux_size3_23_sram[0:1]),
		.mem_outb(clk_mux_size3_23_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_112 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[99:100]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[99:100]),
		.mem_out(clk_mux_size3_24_sram[0:1]),
		.mem_outb(clk_mux_size3_24_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_114 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[101:102]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[101:102]),
		.mem_out(clk_mux_size3_25_sram[0:1]),
		.mem_outb(clk_mux_size3_25_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_116 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[103:104]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[103:104]),
		.mem_out(clk_mux_size3_26_sram[0:1]),
		.mem_outb(clk_mux_size3_26_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_118 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[105:106]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[105:106]),
		.mem_out(clk_mux_size3_27_sram[0:1]),
		.mem_outb(clk_mux_size3_27_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_120 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[107:108]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[107:108]),
		.mem_out(clk_mux_size3_28_sram[0:1]),
		.mem_outb(clk_mux_size3_28_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_122 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[109:110]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[109:110]),
		.mem_out(clk_mux_size3_29_sram[0:1]),
		.mem_outb(clk_mux_size3_29_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_124 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[111:112]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[111:112]),
		.mem_out(clk_mux_size3_30_sram[0:1]),
		.mem_outb(clk_mux_size3_30_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_126 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[113:114]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[113:114]),
		.mem_out(clk_mux_size3_31_sram[0:1]),
		.mem_outb(clk_mux_size3_31_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_65 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[167:168]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[167:168]),
		.mem_out(clk_mux_size3_32_sram[0:1]),
		.mem_outb(clk_mux_size3_32_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_67 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[169:170]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[169:170]),
		.mem_out(clk_mux_size3_33_sram[0:1]),
		.mem_outb(clk_mux_size3_33_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_69 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[171:172]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[171:172]),
		.mem_out(clk_mux_size3_34_sram[0:1]),
		.mem_outb(clk_mux_size3_34_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_71 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[173:174]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[173:174]),
		.mem_out(clk_mux_size3_35_sram[0:1]),
		.mem_outb(clk_mux_size3_35_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_73 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[175:176]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[175:176]),
		.mem_out(clk_mux_size3_36_sram[0:1]),
		.mem_outb(clk_mux_size3_36_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_75 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[177:178]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[177:178]),
		.mem_out(clk_mux_size3_37_sram[0:1]),
		.mem_outb(clk_mux_size3_37_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_77 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[179:180]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[179:180]),
		.mem_out(clk_mux_size3_38_sram[0:1]),
		.mem_outb(clk_mux_size3_38_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_79 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[181:182]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[181:182]),
		.mem_out(clk_mux_size3_39_sram[0:1]),
		.mem_outb(clk_mux_size3_39_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_81 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[183:184]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[183:184]),
		.mem_out(clk_mux_size3_40_sram[0:1]),
		.mem_outb(clk_mux_size3_40_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_83 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[185:186]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[185:186]),
		.mem_out(clk_mux_size3_41_sram[0:1]),
		.mem_outb(clk_mux_size3_41_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_85 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[187:188]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[187:188]),
		.mem_out(clk_mux_size3_42_sram[0:1]),
		.mem_outb(clk_mux_size3_42_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_87 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[189:190]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[189:190]),
		.mem_out(clk_mux_size3_43_sram[0:1]),
		.mem_outb(clk_mux_size3_43_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_89 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[191:192]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[191:192]),
		.mem_out(clk_mux_size3_44_sram[0:1]),
		.mem_outb(clk_mux_size3_44_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_91 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[193:194]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[193:194]),
		.mem_out(clk_mux_size3_45_sram[0:1]),
		.mem_outb(clk_mux_size3_45_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_93 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[195:196]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[195:196]),
		.mem_out(clk_mux_size3_46_sram[0:1]),
		.mem_outb(clk_mux_size3_46_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_95 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[197:198]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[197:198]),
		.mem_out(clk_mux_size3_47_sram[0:1]),
		.mem_outb(clk_mux_size3_47_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_97 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[199:200]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[199:200]),
		.mem_out(clk_mux_size3_48_sram[0:1]),
		.mem_outb(clk_mux_size3_48_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_99 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[201:202]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[201:202]),
		.mem_out(clk_mux_size3_49_sram[0:1]),
		.mem_outb(clk_mux_size3_49_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_101 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[203:204]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[203:204]),
		.mem_out(clk_mux_size3_50_sram[0:1]),
		.mem_outb(clk_mux_size3_50_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_103 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[205:206]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[205:206]),
		.mem_out(clk_mux_size3_51_sram[0:1]),
		.mem_outb(clk_mux_size3_51_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_105 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[207:208]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[207:208]),
		.mem_out(clk_mux_size3_52_sram[0:1]),
		.mem_outb(clk_mux_size3_52_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_107 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[209:210]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[209:210]),
		.mem_out(clk_mux_size3_53_sram[0:1]),
		.mem_outb(clk_mux_size3_53_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_109 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[211:212]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[211:212]),
		.mem_out(clk_mux_size3_54_sram[0:1]),
		.mem_outb(clk_mux_size3_54_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_111 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[213:214]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[213:214]),
		.mem_out(clk_mux_size3_55_sram[0:1]),
		.mem_outb(clk_mux_size3_55_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_113 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[215:216]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[215:216]),
		.mem_out(clk_mux_size3_56_sram[0:1]),
		.mem_outb(clk_mux_size3_56_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_115 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[217:218]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[217:218]),
		.mem_out(clk_mux_size3_57_sram[0:1]),
		.mem_outb(clk_mux_size3_57_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_117 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[219:220]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[219:220]),
		.mem_out(clk_mux_size3_58_sram[0:1]),
		.mem_outb(clk_mux_size3_58_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_119 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[221:222]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[221:222]),
		.mem_out(clk_mux_size3_59_sram[0:1]),
		.mem_outb(clk_mux_size3_59_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_121 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[223:224]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[223:224]),
		.mem_out(clk_mux_size3_60_sram[0:1]),
		.mem_outb(clk_mux_size3_60_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_123 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[225:226]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[225:226]),
		.mem_out(clk_mux_size3_61_sram[0:1]),
		.mem_outb(clk_mux_size3_61_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_125 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[227:228]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[227:228]),
		.mem_out(clk_mux_size3_62_sram[0:1]),
		.mem_outb(clk_mux_size3_62_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_127 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[229:230]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[229:230]),
		.mem_out(clk_mux_size3_63_sram[0:1]),
		.mem_outb(clk_mux_size3_63_sram_inv[0:1]));

	sb_mux_size5 mux_left_track_25 (
		.in({chany_top_in[24], chany_bottom_in[23:24], left_top_grid_bottom_width_0_height_0_subtile_0__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_match1_o_0_}),
		.sram(sb_mux_size5_0_sram[0:2]),
		.sram_inv(sb_mux_size5_0_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	sb_mux_size5 mux_left_track_27 (
		.in({chany_top_in[25], chany_bottom_in[25], chany_bottom_in[27], left_top_grid_bottom_width_0_height_0_subtile_1__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_zero_o_0_}),
		.sram(sb_mux_size5_1_sram[0:2]),
		.sram_inv(sb_mux_size5_1_sram_inv[0:2]),
		.out(chanx_left_out[13]));

	sb_mux_size5 mux_left_track_29 (
		.in({chany_top_in[26], chany_bottom_in[26], chany_bottom_in[31], left_top_grid_bottom_width_0_height_0_subtile_2__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_match1_o_0_}),
		.sram(sb_mux_size5_2_sram[0:2]),
		.sram_inv(sb_mux_size5_2_sram_inv[0:2]),
		.out(chanx_left_out[14]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_25 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[271:273]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[271:273]),
		.mem_out(sb_mux_size5_0_sram[0:2]),
		.mem_outb(sb_mux_size5_0_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_27 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[274:276]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[274:276]),
		.mem_out(sb_mux_size5_1_sram[0:2]),
		.mem_outb(sb_mux_size5_1_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_29 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[277:279]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[277:279]),
		.mem_out(sb_mux_size5_2_sram[0:2]),
		.mem_outb(sb_mux_size5_2_sram_inv[0:2]));

	sb_mux_size4 mux_left_track_31 (
		.in({chany_top_in[28], chany_bottom_in[28], left_top_grid_bottom_width_0_height_0_subtile_3__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_zero_o_0_}),
		.sram(sb_mux_size4_0_sram[0:2]),
		.sram_inv(sb_mux_size4_0_sram_inv[0:2]),
		.out(chanx_left_out[15]));

	sb_mux_size4 mux_left_track_33 (
		.in({chany_top_in[29], chany_bottom_in[29], left_top_grid_bottom_width_0_height_0_subtile_4__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_match1_o_0_}),
		.sram(sb_mux_size4_1_sram[0:2]),
		.sram_inv(sb_mux_size4_1_sram_inv[0:2]),
		.out(chanx_left_out[16]));

	sb_mux_size4 mux_left_track_35 (
		.in({chany_top_in[30], chany_bottom_in[30], left_top_grid_bottom_width_0_height_0_subtile_5__pin_a2f_o_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_zero_o_0_}),
		.sram(sb_mux_size4_2_sram[0:2]),
		.sram_inv(sb_mux_size4_2_sram_inv[0:2]),
		.out(chanx_left_out[17]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_left_track_31 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[280:282]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[280:282]),
		.mem_out(sb_mux_size4_0_sram[0:2]),
		.mem_outb(sb_mux_size4_0_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_left_track_33 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[283:285]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[283:285]),
		.mem_out(sb_mux_size4_1_sram[0:2]),
		.mem_outb(sb_mux_size4_1_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_left_track_35 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[286:288]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[286:288]),
		.mem_out(sb_mux_size4_2_sram[0:2]),
		.mem_outb(sb_mux_size4_2_sram_inv[0:2]));

	sb_mux_size2 mux_left_track_39 (
		.in({chany_top_in[31], left_top_grid_bottom_width_0_height_0_subtile_7__pin_a2f_o_0_}),
		.sram(sb_mux_size2_0_sram[0:1]),
		.sram_inv(sb_mux_size2_0_sram_inv[0:1]),
		.out(chanx_left_out[19]));

	sb_mux_size2 mux_left_track_41 (
		.in({chany_top_in[27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_12_}),
		.sram(sb_mux_size2_1_sram[0:1]),
		.sram_inv(sb_mux_size2_1_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	sb_mux_size2 mux_left_track_43 (
		.in({chany_top_in[23], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_13_}),
		.sram(sb_mux_size2_2_sram[0:1]),
		.sram_inv(sb_mux_size2_2_sram_inv[0:1]),
		.out(chanx_left_out[21]));

	sb_mux_size2 mux_left_track_45 (
		.in({chany_top_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_14_}),
		.sram(sb_mux_size2_3_sram[0:1]),
		.sram_inv(sb_mux_size2_3_sram_inv[0:1]),
		.out(chanx_left_out[22]));

	sb_mux_size2 mux_left_track_47 (
		.in({chany_top_in[15], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_15_}),
		.sram(sb_mux_size2_4_sram[0:1]),
		.sram_inv(sb_mux_size2_4_sram_inv[0:1]),
		.out(chanx_left_out[23]));

	sb_mux_size2 mux_left_track_49 (
		.in({chany_top_in[11], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_16_}),
		.sram(sb_mux_size2_5_sram[0:1]),
		.sram_inv(sb_mux_size2_5_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	sb_mux_size2 mux_left_track_51 (
		.in({chany_top_in[9], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_17_}),
		.sram(sb_mux_size2_6_sram[0:1]),
		.sram_inv(sb_mux_size2_6_sram_inv[0:1]),
		.out(chanx_left_out[25]));

	sb_mux_size2 mux_left_track_53 (
		.in({chany_top_in[7], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_18_}),
		.sram(sb_mux_size2_7_sram[0:1]),
		.sram_inv(sb_mux_size2_7_sram_inv[0:1]),
		.out(chanx_left_out[26]));

	sb_mux_size2 mux_left_track_55 (
		.in({chany_top_in[5], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_19_}),
		.sram(sb_mux_size2_8_sram[0:1]),
		.sram_inv(sb_mux_size2_8_sram_inv[0:1]),
		.out(chanx_left_out[27]));

	sb_mux_size2 mux_left_track_57 (
		.in({chany_top_in[4], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_20_}),
		.sram(sb_mux_size2_9_sram[0:1]),
		.sram_inv(sb_mux_size2_9_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	sb_mux_size2 mux_left_track_59 (
		.in({chany_top_in[3], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_21_}),
		.sram(sb_mux_size2_10_sram[0:1]),
		.sram_inv(sb_mux_size2_10_sram_inv[0:1]),
		.out(chanx_left_out[29]));

	sb_mux_size2 mux_left_track_61 (
		.in({chany_top_in[2], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_22_}),
		.sram(sb_mux_size2_11_sram[0:1]),
		.sram_inv(sb_mux_size2_11_sram_inv[0:1]),
		.out(chanx_left_out[30]));

	sb_mux_size2 mux_left_track_63 (
		.in({chany_top_in[1], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_23_}),
		.sram(sb_mux_size2_12_sram[0:1]),
		.sram_inv(sb_mux_size2_12_sram_inv[0:1]),
		.out(chanx_left_out[31]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_39 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[289:290]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[289:290]),
		.mem_out(sb_mux_size2_0_sram[0:1]),
		.mem_outb(sb_mux_size2_0_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_41 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[291:292]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[291:292]),
		.mem_out(sb_mux_size2_1_sram[0:1]),
		.mem_outb(sb_mux_size2_1_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_43 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[293:294]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[293:294]),
		.mem_out(sb_mux_size2_2_sram[0:1]),
		.mem_outb(sb_mux_size2_2_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_45 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[295:296]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[295:296]),
		.mem_out(sb_mux_size2_3_sram[0:1]),
		.mem_outb(sb_mux_size2_3_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_47 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[297:298]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[297:298]),
		.mem_out(sb_mux_size2_4_sram[0:1]),
		.mem_outb(sb_mux_size2_4_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_49 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[299:300]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[299:300]),
		.mem_out(sb_mux_size2_5_sram[0:1]),
		.mem_outb(sb_mux_size2_5_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_51 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[301:302]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[301:302]),
		.mem_out(sb_mux_size2_6_sram[0:1]),
		.mem_outb(sb_mux_size2_6_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_53 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[303:304]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[303:304]),
		.mem_out(sb_mux_size2_7_sram[0:1]),
		.mem_outb(sb_mux_size2_7_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_55 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[305:306]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[305:306]),
		.mem_out(sb_mux_size2_8_sram[0:1]),
		.mem_outb(sb_mux_size2_8_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_57 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[307:308]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[307:308]),
		.mem_out(sb_mux_size2_9_sram[0:1]),
		.mem_outb(sb_mux_size2_9_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_59 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[309:310]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[309:310]),
		.mem_out(sb_mux_size2_10_sram[0:1]),
		.mem_outb(sb_mux_size2_10_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_61 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[311:312]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[311:312]),
		.mem_out(sb_mux_size2_11_sram[0:1]),
		.mem_outb(sb_mux_size2_11_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_left_track_63 (
		.feedthrough_mem_in(sb_12__config_group_mem_size315_0_mem_out[313:314]),
		.feedthrough_mem_inb(sb_12__config_group_mem_size315_0_mem_outb[313:314]),
		.mem_out(sb_mux_size2_12_sram[0:1]),
		.mem_outb(sb_mux_size2_12_sram_inv[0:1]));

	sb_12__config_group_mem_size315 sb_12__config_group_mem_size315 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.mem_out(sb_12__config_group_mem_size315_0_mem_out[0:314]),
		.mem_outb(sb_12__config_group_mem_size315_0_mem_outb[0:314]),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for sb_12_ -----



