//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Memories used in FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for cb_mux_size8_mem -----
module cb_mux_size8_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for cb_mux_size8_mem -----




// ----- Verilog module for cb_mux_size8_feedthrough_mem -----
module cb_mux_size8_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for cb_mux_size8_feedthrough_mem -----




// ----- Verilog module for cb_mux_size48_mem -----
module cb_mux_size48_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:5] mem_out;
//----- OUTPUT PORTS -----
output [0:5] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

endmodule
// ----- END Verilog module for cb_mux_size48_mem -----




// ----- Verilog module for cb_mux_size48_feedthrough_mem -----
module cb_mux_size48_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:5] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:5] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:5] mem_out;
//----- OUTPUT PORTS -----
output [0:5] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for cb_mux_size48_feedthrough_mem -----




// ----- Verilog module for cb_mux_size16_mem -----
module cb_mux_size16_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

endmodule
// ----- END Verilog module for cb_mux_size16_mem -----




// ----- Verilog module for cb_mux_size16_feedthrough_mem -----
module cb_mux_size16_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for cb_mux_size16_feedthrough_mem -----




// ----- Verilog module for cb_mux_size56_mem -----
module cb_mux_size56_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:5] mem_out;
//----- OUTPUT PORTS -----
output [0:5] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

endmodule
// ----- END Verilog module for cb_mux_size56_mem -----




// ----- Verilog module for cb_mux_size56_feedthrough_mem -----
module cb_mux_size56_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:5] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:5] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:5] mem_out;
//----- OUTPUT PORTS -----
output [0:5] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for cb_mux_size56_feedthrough_mem -----




// ----- Verilog module for cb_mux_size26_mem -----
module cb_mux_size26_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

endmodule
// ----- END Verilog module for cb_mux_size26_mem -----




// ----- Verilog module for cb_mux_size26_feedthrough_mem -----
module cb_mux_size26_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for cb_mux_size26_feedthrough_mem -----




// ----- Verilog module for cb_mux_size76_mem -----
module cb_mux_size76_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(EFPGA_CCFF_5_Q),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

	EFPGA_CCFF EFPGA_CCFF_6_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_5_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[6]),
		.CFGQ(mem_out[6]));

endmodule
// ----- END Verilog module for cb_mux_size76_mem -----




// ----- Verilog module for cb_mux_size76_feedthrough_mem -----
module cb_mux_size76_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[6] = feedthrough_mem_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[6] = feedthrough_mem_inb[6];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for cb_mux_size76_feedthrough_mem -----




// ----- Verilog module for sb_mux_size6_mem -----
module sb_mux_size6_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

endmodule
// ----- END Verilog module for sb_mux_size6_mem -----




// ----- Verilog module for sb_mux_size6_feedthrough_mem -----
module sb_mux_size6_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size6_feedthrough_mem -----




// ----- Verilog module for sb_mux_size5_mem -----
module sb_mux_size5_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

endmodule
// ----- END Verilog module for sb_mux_size5_mem -----




// ----- Verilog module for sb_mux_size5_feedthrough_mem -----
module sb_mux_size5_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size5_feedthrough_mem -----




// ----- Verilog module for sb_mux_size4_mem -----
module sb_mux_size4_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

endmodule
// ----- END Verilog module for sb_mux_size4_mem -----




// ----- Verilog module for sb_mux_size4_feedthrough_mem -----
module sb_mux_size4_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size4_feedthrough_mem -----




// ----- Verilog module for sb_mux_size11_mem -----
module sb_mux_size11_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for sb_mux_size11_mem -----




// ----- Verilog module for sb_mux_size11_feedthrough_mem -----
module sb_mux_size11_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size11_feedthrough_mem -----




// ----- Verilog module for sb_mux_size9_mem -----
module sb_mux_size9_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for sb_mux_size9_mem -----




// ----- Verilog module for sb_mux_size9_feedthrough_mem -----
module sb_mux_size9_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size9_feedthrough_mem -----




// ----- Verilog module for sb_mux_size7_mem -----
module sb_mux_size7_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

endmodule
// ----- END Verilog module for sb_mux_size7_mem -----




// ----- Verilog module for sb_mux_size7_feedthrough_mem -----
module sb_mux_size7_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:2] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:2] mem_out;
//----- OUTPUT PORTS -----
output [0:2] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size7_feedthrough_mem -----




// ----- Verilog module for sb_mux_size8_mem -----
module sb_mux_size8_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for sb_mux_size8_mem -----




// ----- Verilog module for sb_mux_size8_feedthrough_mem -----
module sb_mux_size8_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size8_feedthrough_mem -----




// ----- Verilog module for sb_mux_size10_mem -----
module sb_mux_size10_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for sb_mux_size10_mem -----




// ----- Verilog module for sb_mux_size10_feedthrough_mem -----
module sb_mux_size10_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size10_feedthrough_mem -----




// ----- Verilog module for sb_mux_size17_mem -----
module sb_mux_size17_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

endmodule
// ----- END Verilog module for sb_mux_size17_mem -----




// ----- Verilog module for sb_mux_size17_feedthrough_mem -----
module sb_mux_size17_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size17_feedthrough_mem -----




// ----- Verilog module for sb_mux_size13_mem -----
module sb_mux_size13_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for sb_mux_size13_mem -----




// ----- Verilog module for sb_mux_size13_feedthrough_mem -----
module sb_mux_size13_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size13_feedthrough_mem -----




// ----- Verilog module for sb_mux_size15_mem -----
module sb_mux_size15_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for sb_mux_size15_mem -----




// ----- Verilog module for sb_mux_size15_feedthrough_mem -----
module sb_mux_size15_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size15_feedthrough_mem -----




// ----- Verilog module for sb_mux_size23_mem -----
module sb_mux_size23_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

endmodule
// ----- END Verilog module for sb_mux_size23_mem -----




// ----- Verilog module for sb_mux_size23_feedthrough_mem -----
module sb_mux_size23_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size23_feedthrough_mem -----




// ----- Verilog module for sb_mux_size21_mem -----
module sb_mux_size21_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

endmodule
// ----- END Verilog module for sb_mux_size21_mem -----




// ----- Verilog module for sb_mux_size21_feedthrough_mem -----
module sb_mux_size21_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size21_feedthrough_mem -----




// ----- Verilog module for sb_mux_size3_mem -----
module sb_mux_size3_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

endmodule
// ----- END Verilog module for sb_mux_size3_mem -----




// ----- Verilog module for sb_mux_size3_feedthrough_mem -----
module sb_mux_size3_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size3_feedthrough_mem -----




// ----- Verilog module for sb_mux_size2_mem -----
module sb_mux_size2_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

endmodule
// ----- END Verilog module for sb_mux_size2_mem -----




// ----- Verilog module for sb_mux_size2_feedthrough_mem -----
module sb_mux_size2_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size2_feedthrough_mem -----




// ----- Verilog module for sb_mux_size12_mem -----
module sb_mux_size12_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for sb_mux_size12_mem -----




// ----- Verilog module for sb_mux_size12_feedthrough_mem -----
module sb_mux_size12_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size12_feedthrough_mem -----




// ----- Verilog module for sb_mux_size19_mem -----
module sb_mux_size19_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

endmodule
// ----- END Verilog module for sb_mux_size19_mem -----




// ----- Verilog module for sb_mux_size19_feedthrough_mem -----
module sb_mux_size19_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for sb_mux_size19_feedthrough_mem -----




// ----- Verilog module for clk_mux_size3_mem -----
module clk_mux_size3_mem(config_enable,
                         prog_reset,
                         prog_clk,
                         ccff_head,
                         ccff_tail,
                         mem_out,
                         mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

endmodule
// ----- END Verilog module for clk_mux_size3_mem -----




// ----- Verilog module for clk_mux_size3_feedthrough_mem -----
module clk_mux_size3_feedthrough_mem(feedthrough_mem_in,
                                     feedthrough_mem_inb,
                                     mem_out,
                                     mem_outb);
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for clk_mux_size3_feedthrough_mem -----




// ----- Verilog module for pb_mux_highload_size2_mem -----
module pb_mux_highload_size2_mem(config_enable,
                                 prog_reset,
                                 prog_clk,
                                 ccff_head,
                                 ccff_tail,
                                 mem_out,
                                 mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:0] mem_out;
//----- OUTPUT PORTS -----
output [0:0] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(ccff_tail),
		.CFGQN(mem_outb),
		.CFGQ(mem_out));

endmodule
// ----- END Verilog module for pb_mux_highload_size2_mem -----




// ----- Verilog module for pb_mux_highload_size2_feedthrough_mem -----
module pb_mux_highload_size2_feedthrough_mem(feedthrough_mem_in,
                                             feedthrough_mem_inb,
                                             mem_out,
                                             mem_outb);
//----- INPUT PORTS -----
input [0:0] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:0] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:0] mem_out;
//----- OUTPUT PORTS -----
output [0:0] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for pb_mux_highload_size2_feedthrough_mem -----




// ----- Verilog module for pb_mux_highload_size3_mem -----
module pb_mux_highload_size3_mem(config_enable,
                                 prog_reset,
                                 prog_clk,
                                 ccff_head,
                                 ccff_tail,
                                 mem_out,
                                 mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

endmodule
// ----- END Verilog module for pb_mux_highload_size3_mem -----




// ----- Verilog module for pb_mux_highload_size3_feedthrough_mem -----
module pb_mux_highload_size3_feedthrough_mem(feedthrough_mem_in,
                                             feedthrough_mem_inb,
                                             mem_out,
                                             mem_outb);
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for pb_mux_highload_size3_feedthrough_mem -----




// ----- Verilog module for pb_mux_no_const_input_size2_mem -----
module pb_mux_no_const_input_size2_mem(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       ccff_tail,
                                       mem_out,
                                       mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:0] mem_out;
//----- OUTPUT PORTS -----
output [0:0] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(ccff_tail),
		.CFGQN(mem_outb),
		.CFGQ(mem_out));

endmodule
// ----- END Verilog module for pb_mux_no_const_input_size2_mem -----




// ----- Verilog module for pb_mux_no_const_input_size2_feedthrough_mem -----
module pb_mux_no_const_input_size2_feedthrough_mem(feedthrough_mem_in,
                                                   feedthrough_mem_inb,
                                                   mem_out,
                                                   mem_outb);
//----- INPUT PORTS -----
input [0:0] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:0] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:0] mem_out;
//----- OUTPUT PORTS -----
output [0:0] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for pb_mux_no_const_input_size2_feedthrough_mem -----




// ----- Verilog module for pb_mux_size2_mem -----
module pb_mux_size2_mem(config_enable,
                        prog_reset,
                        prog_clk,
                        ccff_head,
                        ccff_tail,
                        mem_out,
                        mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

endmodule
// ----- END Verilog module for pb_mux_size2_mem -----




// ----- Verilog module for pb_mux_size2_feedthrough_mem -----
module pb_mux_size2_feedthrough_mem(feedthrough_mem_in,
                                    feedthrough_mem_inb,
                                    mem_out,
                                    mem_outb);
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:1] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:1] mem_out;
//----- OUTPUT PORTS -----
output [0:1] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for pb_mux_size2_feedthrough_mem -----




// ----- Verilog module for mmff_wrapper_EFPGA_CCFF_mem -----
module mmff_wrapper_EFPGA_CCFF_mem(config_enable,
                                   prog_reset,
                                   prog_clk,
                                   ccff_head,
                                   ccff_tail,
                                   mem_out,
                                   mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

endmodule
// ----- END Verilog module for mmff_wrapper_EFPGA_CCFF_mem -----




// ----- Verilog module for mmff_wrapper_feedthrough_EFPGA_CCFF_mem -----
module mmff_wrapper_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                               feedthrough_mem_inb,
                                               mem_out,
                                               mem_outb);
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:3] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:3] mem_out;
//----- OUTPUT PORTS -----
output [0:3] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for mmff_wrapper_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for mmffisc2_wrapper_EFPGA_CCFF_mem -----
module mmffisc2_wrapper_EFPGA_CCFF_mem(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       ccff_tail,
                                       mem_out,
                                       mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(EFPGA_CCFF_5_Q),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

	EFPGA_CCFF EFPGA_CCFF_6_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_5_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[6]),
		.CFGQ(mem_out[6]));

endmodule
// ----- END Verilog module for mmffisc2_wrapper_EFPGA_CCFF_mem -----




// ----- Verilog module for mmffisc2_wrapper_feedthrough_EFPGA_CCFF_mem -----
module mmffisc2_wrapper_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                                   feedthrough_mem_inb,
                                                   mem_out,
                                                   mem_outb);
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[6] = feedthrough_mem_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[6] = feedthrough_mem_inb[6];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for mmffisc2_wrapper_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for mmffosc2_wrapper_EFPGA_CCFF_mem -----
module mmffosc2_wrapper_EFPGA_CCFF_mem(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       ccff_tail,
                                       mem_out,
                                       mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(EFPGA_CCFF_5_Q),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

	EFPGA_CCFF EFPGA_CCFF_6_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_5_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[6]),
		.CFGQ(mem_out[6]));

endmodule
// ----- END Verilog module for mmffosc2_wrapper_EFPGA_CCFF_mem -----




// ----- Verilog module for mmffosc2_wrapper_feedthrough_EFPGA_CCFF_mem -----
module mmffosc2_wrapper_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                                   feedthrough_mem_inb,
                                                   mem_out,
                                                   mem_outb);
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[6] = feedthrough_mem_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[6] = feedthrough_mem_inb[6];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for mmffosc2_wrapper_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for mmffosc2cko_wrapper_EFPGA_CCFF_mem -----
module mmffosc2cko_wrapper_EFPGA_CCFF_mem(config_enable,
                                          prog_reset,
                                          prog_clk,
                                          ccff_head,
                                          ccff_tail,
                                          mem_out,
                                          mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(EFPGA_CCFF_5_Q),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

	EFPGA_CCFF EFPGA_CCFF_6_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_5_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[6]),
		.CFGQ(mem_out[6]));

endmodule
// ----- END Verilog module for mmffosc2cko_wrapper_EFPGA_CCFF_mem -----




// ----- Verilog module for mmffosc2cko_wrapper_feedthrough_EFPGA_CCFF_mem -----
module mmffosc2cko_wrapper_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                                      feedthrough_mem_inb,
                                                      mem_out,
                                                      mem_outb);
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:6] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:6] mem_out;
//----- OUTPUT PORTS -----
output [0:6] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[6] = feedthrough_mem_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[6] = feedthrough_mem_inb[6];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for mmffosc2cko_wrapper_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for frac_lut5_arith_EFPGA_CCFF_mem -----
module frac_lut5_arith_EFPGA_CCFF_mem(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      ccff_tail,
                                      mem_out,
                                      mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:32] mem_out;
//----- OUTPUT PORTS -----
output [0:32] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(EFPGA_CCFF_5_Q),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

	EFPGA_CCFF EFPGA_CCFF_6_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_5_Q),
		.Q(EFPGA_CCFF_6_Q),
		.CFGQN(mem_outb[6]),
		.CFGQ(mem_out[6]));

	EFPGA_CCFF EFPGA_CCFF_7_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_6_Q),
		.Q(EFPGA_CCFF_7_Q),
		.CFGQN(mem_outb[7]),
		.CFGQ(mem_out[7]));

	EFPGA_CCFF EFPGA_CCFF_8_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_7_Q),
		.Q(EFPGA_CCFF_8_Q),
		.CFGQN(mem_outb[8]),
		.CFGQ(mem_out[8]));

	EFPGA_CCFF EFPGA_CCFF_9_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_8_Q),
		.Q(EFPGA_CCFF_9_Q),
		.CFGQN(mem_outb[9]),
		.CFGQ(mem_out[9]));

	EFPGA_CCFF EFPGA_CCFF_10_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_9_Q),
		.Q(EFPGA_CCFF_10_Q),
		.CFGQN(mem_outb[10]),
		.CFGQ(mem_out[10]));

	EFPGA_CCFF EFPGA_CCFF_11_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_10_Q),
		.Q(EFPGA_CCFF_11_Q),
		.CFGQN(mem_outb[11]),
		.CFGQ(mem_out[11]));

	EFPGA_CCFF EFPGA_CCFF_12_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_11_Q),
		.Q(EFPGA_CCFF_12_Q),
		.CFGQN(mem_outb[12]),
		.CFGQ(mem_out[12]));

	EFPGA_CCFF EFPGA_CCFF_13_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_12_Q),
		.Q(EFPGA_CCFF_13_Q),
		.CFGQN(mem_outb[13]),
		.CFGQ(mem_out[13]));

	EFPGA_CCFF EFPGA_CCFF_14_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_13_Q),
		.Q(EFPGA_CCFF_14_Q),
		.CFGQN(mem_outb[14]),
		.CFGQ(mem_out[14]));

	EFPGA_CCFF EFPGA_CCFF_15_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_14_Q),
		.Q(EFPGA_CCFF_15_Q),
		.CFGQN(mem_outb[15]),
		.CFGQ(mem_out[15]));

	EFPGA_CCFF EFPGA_CCFF_16_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_15_Q),
		.Q(EFPGA_CCFF_16_Q),
		.CFGQN(mem_outb[16]),
		.CFGQ(mem_out[16]));

	EFPGA_CCFF EFPGA_CCFF_17_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_16_Q),
		.Q(EFPGA_CCFF_17_Q),
		.CFGQN(mem_outb[17]),
		.CFGQ(mem_out[17]));

	EFPGA_CCFF EFPGA_CCFF_18_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_17_Q),
		.Q(EFPGA_CCFF_18_Q),
		.CFGQN(mem_outb[18]),
		.CFGQ(mem_out[18]));

	EFPGA_CCFF EFPGA_CCFF_19_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_18_Q),
		.Q(EFPGA_CCFF_19_Q),
		.CFGQN(mem_outb[19]),
		.CFGQ(mem_out[19]));

	EFPGA_CCFF EFPGA_CCFF_20_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_19_Q),
		.Q(EFPGA_CCFF_20_Q),
		.CFGQN(mem_outb[20]),
		.CFGQ(mem_out[20]));

	EFPGA_CCFF EFPGA_CCFF_21_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_20_Q),
		.Q(EFPGA_CCFF_21_Q),
		.CFGQN(mem_outb[21]),
		.CFGQ(mem_out[21]));

	EFPGA_CCFF EFPGA_CCFF_22_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_21_Q),
		.Q(EFPGA_CCFF_22_Q),
		.CFGQN(mem_outb[22]),
		.CFGQ(mem_out[22]));

	EFPGA_CCFF EFPGA_CCFF_23_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_22_Q),
		.Q(EFPGA_CCFF_23_Q),
		.CFGQN(mem_outb[23]),
		.CFGQ(mem_out[23]));

	EFPGA_CCFF EFPGA_CCFF_24_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_23_Q),
		.Q(EFPGA_CCFF_24_Q),
		.CFGQN(mem_outb[24]),
		.CFGQ(mem_out[24]));

	EFPGA_CCFF EFPGA_CCFF_25_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_24_Q),
		.Q(EFPGA_CCFF_25_Q),
		.CFGQN(mem_outb[25]),
		.CFGQ(mem_out[25]));

	EFPGA_CCFF EFPGA_CCFF_26_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_25_Q),
		.Q(EFPGA_CCFF_26_Q),
		.CFGQN(mem_outb[26]),
		.CFGQ(mem_out[26]));

	EFPGA_CCFF EFPGA_CCFF_27_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_26_Q),
		.Q(EFPGA_CCFF_27_Q),
		.CFGQN(mem_outb[27]),
		.CFGQ(mem_out[27]));

	EFPGA_CCFF EFPGA_CCFF_28_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_27_Q),
		.Q(EFPGA_CCFF_28_Q),
		.CFGQN(mem_outb[28]),
		.CFGQ(mem_out[28]));

	EFPGA_CCFF EFPGA_CCFF_29_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_28_Q),
		.Q(EFPGA_CCFF_29_Q),
		.CFGQN(mem_outb[29]),
		.CFGQ(mem_out[29]));

	EFPGA_CCFF EFPGA_CCFF_30_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_29_Q),
		.Q(EFPGA_CCFF_30_Q),
		.CFGQN(mem_outb[30]),
		.CFGQ(mem_out[30]));

	EFPGA_CCFF EFPGA_CCFF_31_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_30_Q),
		.Q(EFPGA_CCFF_31_Q),
		.CFGQN(mem_outb[31]),
		.CFGQ(mem_out[31]));

	EFPGA_CCFF EFPGA_CCFF_32_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_31_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[32]),
		.CFGQ(mem_out[32]));

endmodule
// ----- END Verilog module for frac_lut5_arith_EFPGA_CCFF_mem -----




// ----- Verilog module for frac_lut5_arith_feedthrough_EFPGA_CCFF_mem -----
module frac_lut5_arith_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                                  feedthrough_mem_inb,
                                                  mem_out,
                                                  mem_outb);
//----- INPUT PORTS -----
input [0:32] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:32] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:32] mem_out;
//----- OUTPUT PORTS -----
output [0:32] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[6] = feedthrough_mem_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[7] = feedthrough_mem_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[8] = feedthrough_mem_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[9] = feedthrough_mem_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[10] = feedthrough_mem_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[11] = feedthrough_mem_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[12] = feedthrough_mem_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[13] = feedthrough_mem_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[14] = feedthrough_mem_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[15] = feedthrough_mem_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[16] = feedthrough_mem_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[17] = feedthrough_mem_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[18] = feedthrough_mem_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[19] = feedthrough_mem_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[20] = feedthrough_mem_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[21] = feedthrough_mem_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[22] = feedthrough_mem_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[23] = feedthrough_mem_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[24] = feedthrough_mem_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[25] = feedthrough_mem_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[26] = feedthrough_mem_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[27] = feedthrough_mem_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[28] = feedthrough_mem_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[29] = feedthrough_mem_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[30] = feedthrough_mem_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[31] = feedthrough_mem_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[32] = feedthrough_mem_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[6] = feedthrough_mem_inb[6];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[7] = feedthrough_mem_inb[7];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[8] = feedthrough_mem_inb[8];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[9] = feedthrough_mem_inb[9];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[10] = feedthrough_mem_inb[10];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[11] = feedthrough_mem_inb[11];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[12] = feedthrough_mem_inb[12];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[13] = feedthrough_mem_inb[13];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[14] = feedthrough_mem_inb[14];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[15] = feedthrough_mem_inb[15];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[16] = feedthrough_mem_inb[16];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[17] = feedthrough_mem_inb[17];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[18] = feedthrough_mem_inb[18];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[19] = feedthrough_mem_inb[19];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[20] = feedthrough_mem_inb[20];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[21] = feedthrough_mem_inb[21];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[22] = feedthrough_mem_inb[22];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[23] = feedthrough_mem_inb[23];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[24] = feedthrough_mem_inb[24];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[25] = feedthrough_mem_inb[25];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[26] = feedthrough_mem_inb[26];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[27] = feedthrough_mem_inb[27];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[28] = feedthrough_mem_inb[28];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[29] = feedthrough_mem_inb[29];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[30] = feedthrough_mem_inb[30];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[31] = feedthrough_mem_inb[31];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[32] = feedthrough_mem_inb[32];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for frac_lut5_arith_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for pinput_extmode_EFPGA_CCFF_mem -----
module pinput_extmode_EFPGA_CCFF_mem(config_enable,
                                     prog_reset,
                                     prog_clk,
                                     ccff_head,
                                     ccff_tail,
                                     mem_out,
                                     mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:0] mem_out;
//----- OUTPUT PORTS -----
output [0:0] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(ccff_tail),
		.CFGQN(mem_outb),
		.CFGQ(mem_out));

endmodule
// ----- END Verilog module for pinput_extmode_EFPGA_CCFF_mem -----




// ----- Verilog module for pinput_extmode_feedthrough_EFPGA_CCFF_mem -----
module pinput_extmode_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                                 feedthrough_mem_inb,
                                                 mem_out,
                                                 mem_outb);
//----- INPUT PORTS -----
input [0:0] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:0] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:0] mem_out;
//----- OUTPUT PORTS -----
output [0:0] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for pinput_extmode_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for pinput_dchain_extmode_EFPGA_CCFF_mem -----
module pinput_dchain_extmode_EFPGA_CCFF_mem(config_enable,
                                            prog_reset,
                                            prog_clk,
                                            ccff_head,
                                            ccff_tail,
                                            mem_out,
                                            mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

endmodule
// ----- END Verilog module for pinput_dchain_extmode_EFPGA_CCFF_mem -----




// ----- Verilog module for pinput_dchain_extmode_feedthrough_EFPGA_CCFF_mem -----
module pinput_dchain_extmode_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                                        feedthrough_mem_inb,
                                                        mem_out,
                                                        mem_outb);
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:4] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:4] mem_out;
//----- OUTPUT PORTS -----
output [0:4] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for pinput_dchain_extmode_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for pcnt_wrapper_EFPGA_CCFF_mem -----
module pcnt_wrapper_EFPGA_CCFF_mem(config_enable,
                                   prog_reset,
                                   prog_clk,
                                   ccff_head,
                                   ccff_tail,
                                   mem_out,
                                   mem_outb);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;
//----- OUTPUT PORTS -----
output [0:106] mem_out;
//----- OUTPUT PORTS -----
output [0:106] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	EFPGA_CCFF EFPGA_CCFF_0_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(ccff_head),
		.Q(EFPGA_CCFF_0_Q),
		.CFGQN(mem_outb[0]),
		.CFGQ(mem_out[0]));

	EFPGA_CCFF EFPGA_CCFF_1_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_0_Q),
		.Q(EFPGA_CCFF_1_Q),
		.CFGQN(mem_outb[1]),
		.CFGQ(mem_out[1]));

	EFPGA_CCFF EFPGA_CCFF_2_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_1_Q),
		.Q(EFPGA_CCFF_2_Q),
		.CFGQN(mem_outb[2]),
		.CFGQ(mem_out[2]));

	EFPGA_CCFF EFPGA_CCFF_3_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_2_Q),
		.Q(EFPGA_CCFF_3_Q),
		.CFGQN(mem_outb[3]),
		.CFGQ(mem_out[3]));

	EFPGA_CCFF EFPGA_CCFF_4_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_3_Q),
		.Q(EFPGA_CCFF_4_Q),
		.CFGQN(mem_outb[4]),
		.CFGQ(mem_out[4]));

	EFPGA_CCFF EFPGA_CCFF_5_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_4_Q),
		.Q(EFPGA_CCFF_5_Q),
		.CFGQN(mem_outb[5]),
		.CFGQ(mem_out[5]));

	EFPGA_CCFF EFPGA_CCFF_6_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_5_Q),
		.Q(EFPGA_CCFF_6_Q),
		.CFGQN(mem_outb[6]),
		.CFGQ(mem_out[6]));

	EFPGA_CCFF EFPGA_CCFF_7_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_6_Q),
		.Q(EFPGA_CCFF_7_Q),
		.CFGQN(mem_outb[7]),
		.CFGQ(mem_out[7]));

	EFPGA_CCFF EFPGA_CCFF_8_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_7_Q),
		.Q(EFPGA_CCFF_8_Q),
		.CFGQN(mem_outb[8]),
		.CFGQ(mem_out[8]));

	EFPGA_CCFF EFPGA_CCFF_9_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_8_Q),
		.Q(EFPGA_CCFF_9_Q),
		.CFGQN(mem_outb[9]),
		.CFGQ(mem_out[9]));

	EFPGA_CCFF EFPGA_CCFF_10_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_9_Q),
		.Q(EFPGA_CCFF_10_Q),
		.CFGQN(mem_outb[10]),
		.CFGQ(mem_out[10]));

	EFPGA_CCFF EFPGA_CCFF_11_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_10_Q),
		.Q(EFPGA_CCFF_11_Q),
		.CFGQN(mem_outb[11]),
		.CFGQ(mem_out[11]));

	EFPGA_CCFF EFPGA_CCFF_12_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_11_Q),
		.Q(EFPGA_CCFF_12_Q),
		.CFGQN(mem_outb[12]),
		.CFGQ(mem_out[12]));

	EFPGA_CCFF EFPGA_CCFF_13_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_12_Q),
		.Q(EFPGA_CCFF_13_Q),
		.CFGQN(mem_outb[13]),
		.CFGQ(mem_out[13]));

	EFPGA_CCFF EFPGA_CCFF_14_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_13_Q),
		.Q(EFPGA_CCFF_14_Q),
		.CFGQN(mem_outb[14]),
		.CFGQ(mem_out[14]));

	EFPGA_CCFF EFPGA_CCFF_15_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_14_Q),
		.Q(EFPGA_CCFF_15_Q),
		.CFGQN(mem_outb[15]),
		.CFGQ(mem_out[15]));

	EFPGA_CCFF EFPGA_CCFF_16_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_15_Q),
		.Q(EFPGA_CCFF_16_Q),
		.CFGQN(mem_outb[16]),
		.CFGQ(mem_out[16]));

	EFPGA_CCFF EFPGA_CCFF_17_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_16_Q),
		.Q(EFPGA_CCFF_17_Q),
		.CFGQN(mem_outb[17]),
		.CFGQ(mem_out[17]));

	EFPGA_CCFF EFPGA_CCFF_18_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_17_Q),
		.Q(EFPGA_CCFF_18_Q),
		.CFGQN(mem_outb[18]),
		.CFGQ(mem_out[18]));

	EFPGA_CCFF EFPGA_CCFF_19_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_18_Q),
		.Q(EFPGA_CCFF_19_Q),
		.CFGQN(mem_outb[19]),
		.CFGQ(mem_out[19]));

	EFPGA_CCFF EFPGA_CCFF_20_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_19_Q),
		.Q(EFPGA_CCFF_20_Q),
		.CFGQN(mem_outb[20]),
		.CFGQ(mem_out[20]));

	EFPGA_CCFF EFPGA_CCFF_21_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_20_Q),
		.Q(EFPGA_CCFF_21_Q),
		.CFGQN(mem_outb[21]),
		.CFGQ(mem_out[21]));

	EFPGA_CCFF EFPGA_CCFF_22_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_21_Q),
		.Q(EFPGA_CCFF_22_Q),
		.CFGQN(mem_outb[22]),
		.CFGQ(mem_out[22]));

	EFPGA_CCFF EFPGA_CCFF_23_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_22_Q),
		.Q(EFPGA_CCFF_23_Q),
		.CFGQN(mem_outb[23]),
		.CFGQ(mem_out[23]));

	EFPGA_CCFF EFPGA_CCFF_24_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_23_Q),
		.Q(EFPGA_CCFF_24_Q),
		.CFGQN(mem_outb[24]),
		.CFGQ(mem_out[24]));

	EFPGA_CCFF EFPGA_CCFF_25_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_24_Q),
		.Q(EFPGA_CCFF_25_Q),
		.CFGQN(mem_outb[25]),
		.CFGQ(mem_out[25]));

	EFPGA_CCFF EFPGA_CCFF_26_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_25_Q),
		.Q(EFPGA_CCFF_26_Q),
		.CFGQN(mem_outb[26]),
		.CFGQ(mem_out[26]));

	EFPGA_CCFF EFPGA_CCFF_27_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_26_Q),
		.Q(EFPGA_CCFF_27_Q),
		.CFGQN(mem_outb[27]),
		.CFGQ(mem_out[27]));

	EFPGA_CCFF EFPGA_CCFF_28_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_27_Q),
		.Q(EFPGA_CCFF_28_Q),
		.CFGQN(mem_outb[28]),
		.CFGQ(mem_out[28]));

	EFPGA_CCFF EFPGA_CCFF_29_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_28_Q),
		.Q(EFPGA_CCFF_29_Q),
		.CFGQN(mem_outb[29]),
		.CFGQ(mem_out[29]));

	EFPGA_CCFF EFPGA_CCFF_30_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_29_Q),
		.Q(EFPGA_CCFF_30_Q),
		.CFGQN(mem_outb[30]),
		.CFGQ(mem_out[30]));

	EFPGA_CCFF EFPGA_CCFF_31_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_30_Q),
		.Q(EFPGA_CCFF_31_Q),
		.CFGQN(mem_outb[31]),
		.CFGQ(mem_out[31]));

	EFPGA_CCFF EFPGA_CCFF_32_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_31_Q),
		.Q(EFPGA_CCFF_32_Q),
		.CFGQN(mem_outb[32]),
		.CFGQ(mem_out[32]));

	EFPGA_CCFF EFPGA_CCFF_33_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_32_Q),
		.Q(EFPGA_CCFF_33_Q),
		.CFGQN(mem_outb[33]),
		.CFGQ(mem_out[33]));

	EFPGA_CCFF EFPGA_CCFF_34_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_33_Q),
		.Q(EFPGA_CCFF_34_Q),
		.CFGQN(mem_outb[34]),
		.CFGQ(mem_out[34]));

	EFPGA_CCFF EFPGA_CCFF_35_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_34_Q),
		.Q(EFPGA_CCFF_35_Q),
		.CFGQN(mem_outb[35]),
		.CFGQ(mem_out[35]));

	EFPGA_CCFF EFPGA_CCFF_36_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_35_Q),
		.Q(EFPGA_CCFF_36_Q),
		.CFGQN(mem_outb[36]),
		.CFGQ(mem_out[36]));

	EFPGA_CCFF EFPGA_CCFF_37_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_36_Q),
		.Q(EFPGA_CCFF_37_Q),
		.CFGQN(mem_outb[37]),
		.CFGQ(mem_out[37]));

	EFPGA_CCFF EFPGA_CCFF_38_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_37_Q),
		.Q(EFPGA_CCFF_38_Q),
		.CFGQN(mem_outb[38]),
		.CFGQ(mem_out[38]));

	EFPGA_CCFF EFPGA_CCFF_39_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_38_Q),
		.Q(EFPGA_CCFF_39_Q),
		.CFGQN(mem_outb[39]),
		.CFGQ(mem_out[39]));

	EFPGA_CCFF EFPGA_CCFF_40_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_39_Q),
		.Q(EFPGA_CCFF_40_Q),
		.CFGQN(mem_outb[40]),
		.CFGQ(mem_out[40]));

	EFPGA_CCFF EFPGA_CCFF_41_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_40_Q),
		.Q(EFPGA_CCFF_41_Q),
		.CFGQN(mem_outb[41]),
		.CFGQ(mem_out[41]));

	EFPGA_CCFF EFPGA_CCFF_42_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_41_Q),
		.Q(EFPGA_CCFF_42_Q),
		.CFGQN(mem_outb[42]),
		.CFGQ(mem_out[42]));

	EFPGA_CCFF EFPGA_CCFF_43_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_42_Q),
		.Q(EFPGA_CCFF_43_Q),
		.CFGQN(mem_outb[43]),
		.CFGQ(mem_out[43]));

	EFPGA_CCFF EFPGA_CCFF_44_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_43_Q),
		.Q(EFPGA_CCFF_44_Q),
		.CFGQN(mem_outb[44]),
		.CFGQ(mem_out[44]));

	EFPGA_CCFF EFPGA_CCFF_45_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_44_Q),
		.Q(EFPGA_CCFF_45_Q),
		.CFGQN(mem_outb[45]),
		.CFGQ(mem_out[45]));

	EFPGA_CCFF EFPGA_CCFF_46_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_45_Q),
		.Q(EFPGA_CCFF_46_Q),
		.CFGQN(mem_outb[46]),
		.CFGQ(mem_out[46]));

	EFPGA_CCFF EFPGA_CCFF_47_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_46_Q),
		.Q(EFPGA_CCFF_47_Q),
		.CFGQN(mem_outb[47]),
		.CFGQ(mem_out[47]));

	EFPGA_CCFF EFPGA_CCFF_48_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_47_Q),
		.Q(EFPGA_CCFF_48_Q),
		.CFGQN(mem_outb[48]),
		.CFGQ(mem_out[48]));

	EFPGA_CCFF EFPGA_CCFF_49_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_48_Q),
		.Q(EFPGA_CCFF_49_Q),
		.CFGQN(mem_outb[49]),
		.CFGQ(mem_out[49]));

	EFPGA_CCFF EFPGA_CCFF_50_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_49_Q),
		.Q(EFPGA_CCFF_50_Q),
		.CFGQN(mem_outb[50]),
		.CFGQ(mem_out[50]));

	EFPGA_CCFF EFPGA_CCFF_51_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_50_Q),
		.Q(EFPGA_CCFF_51_Q),
		.CFGQN(mem_outb[51]),
		.CFGQ(mem_out[51]));

	EFPGA_CCFF EFPGA_CCFF_52_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_51_Q),
		.Q(EFPGA_CCFF_52_Q),
		.CFGQN(mem_outb[52]),
		.CFGQ(mem_out[52]));

	EFPGA_CCFF EFPGA_CCFF_53_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_52_Q),
		.Q(EFPGA_CCFF_53_Q),
		.CFGQN(mem_outb[53]),
		.CFGQ(mem_out[53]));

	EFPGA_CCFF EFPGA_CCFF_54_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_53_Q),
		.Q(EFPGA_CCFF_54_Q),
		.CFGQN(mem_outb[54]),
		.CFGQ(mem_out[54]));

	EFPGA_CCFF EFPGA_CCFF_55_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_54_Q),
		.Q(EFPGA_CCFF_55_Q),
		.CFGQN(mem_outb[55]),
		.CFGQ(mem_out[55]));

	EFPGA_CCFF EFPGA_CCFF_56_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_55_Q),
		.Q(EFPGA_CCFF_56_Q),
		.CFGQN(mem_outb[56]),
		.CFGQ(mem_out[56]));

	EFPGA_CCFF EFPGA_CCFF_57_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_56_Q),
		.Q(EFPGA_CCFF_57_Q),
		.CFGQN(mem_outb[57]),
		.CFGQ(mem_out[57]));

	EFPGA_CCFF EFPGA_CCFF_58_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_57_Q),
		.Q(EFPGA_CCFF_58_Q),
		.CFGQN(mem_outb[58]),
		.CFGQ(mem_out[58]));

	EFPGA_CCFF EFPGA_CCFF_59_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_58_Q),
		.Q(EFPGA_CCFF_59_Q),
		.CFGQN(mem_outb[59]),
		.CFGQ(mem_out[59]));

	EFPGA_CCFF EFPGA_CCFF_60_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_59_Q),
		.Q(EFPGA_CCFF_60_Q),
		.CFGQN(mem_outb[60]),
		.CFGQ(mem_out[60]));

	EFPGA_CCFF EFPGA_CCFF_61_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_60_Q),
		.Q(EFPGA_CCFF_61_Q),
		.CFGQN(mem_outb[61]),
		.CFGQ(mem_out[61]));

	EFPGA_CCFF EFPGA_CCFF_62_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_61_Q),
		.Q(EFPGA_CCFF_62_Q),
		.CFGQN(mem_outb[62]),
		.CFGQ(mem_out[62]));

	EFPGA_CCFF EFPGA_CCFF_63_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_62_Q),
		.Q(EFPGA_CCFF_63_Q),
		.CFGQN(mem_outb[63]),
		.CFGQ(mem_out[63]));

	EFPGA_CCFF EFPGA_CCFF_64_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_63_Q),
		.Q(EFPGA_CCFF_64_Q),
		.CFGQN(mem_outb[64]),
		.CFGQ(mem_out[64]));

	EFPGA_CCFF EFPGA_CCFF_65_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_64_Q),
		.Q(EFPGA_CCFF_65_Q),
		.CFGQN(mem_outb[65]),
		.CFGQ(mem_out[65]));

	EFPGA_CCFF EFPGA_CCFF_66_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_65_Q),
		.Q(EFPGA_CCFF_66_Q),
		.CFGQN(mem_outb[66]),
		.CFGQ(mem_out[66]));

	EFPGA_CCFF EFPGA_CCFF_67_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_66_Q),
		.Q(EFPGA_CCFF_67_Q),
		.CFGQN(mem_outb[67]),
		.CFGQ(mem_out[67]));

	EFPGA_CCFF EFPGA_CCFF_68_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_67_Q),
		.Q(EFPGA_CCFF_68_Q),
		.CFGQN(mem_outb[68]),
		.CFGQ(mem_out[68]));

	EFPGA_CCFF EFPGA_CCFF_69_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_68_Q),
		.Q(EFPGA_CCFF_69_Q),
		.CFGQN(mem_outb[69]),
		.CFGQ(mem_out[69]));

	EFPGA_CCFF EFPGA_CCFF_70_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_69_Q),
		.Q(EFPGA_CCFF_70_Q),
		.CFGQN(mem_outb[70]),
		.CFGQ(mem_out[70]));

	EFPGA_CCFF EFPGA_CCFF_71_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_70_Q),
		.Q(EFPGA_CCFF_71_Q),
		.CFGQN(mem_outb[71]),
		.CFGQ(mem_out[71]));

	EFPGA_CCFF EFPGA_CCFF_72_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_71_Q),
		.Q(EFPGA_CCFF_72_Q),
		.CFGQN(mem_outb[72]),
		.CFGQ(mem_out[72]));

	EFPGA_CCFF EFPGA_CCFF_73_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_72_Q),
		.Q(EFPGA_CCFF_73_Q),
		.CFGQN(mem_outb[73]),
		.CFGQ(mem_out[73]));

	EFPGA_CCFF EFPGA_CCFF_74_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_73_Q),
		.Q(EFPGA_CCFF_74_Q),
		.CFGQN(mem_outb[74]),
		.CFGQ(mem_out[74]));

	EFPGA_CCFF EFPGA_CCFF_75_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_74_Q),
		.Q(EFPGA_CCFF_75_Q),
		.CFGQN(mem_outb[75]),
		.CFGQ(mem_out[75]));

	EFPGA_CCFF EFPGA_CCFF_76_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_75_Q),
		.Q(EFPGA_CCFF_76_Q),
		.CFGQN(mem_outb[76]),
		.CFGQ(mem_out[76]));

	EFPGA_CCFF EFPGA_CCFF_77_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_76_Q),
		.Q(EFPGA_CCFF_77_Q),
		.CFGQN(mem_outb[77]),
		.CFGQ(mem_out[77]));

	EFPGA_CCFF EFPGA_CCFF_78_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_77_Q),
		.Q(EFPGA_CCFF_78_Q),
		.CFGQN(mem_outb[78]),
		.CFGQ(mem_out[78]));

	EFPGA_CCFF EFPGA_CCFF_79_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_78_Q),
		.Q(EFPGA_CCFF_79_Q),
		.CFGQN(mem_outb[79]),
		.CFGQ(mem_out[79]));

	EFPGA_CCFF EFPGA_CCFF_80_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_79_Q),
		.Q(EFPGA_CCFF_80_Q),
		.CFGQN(mem_outb[80]),
		.CFGQ(mem_out[80]));

	EFPGA_CCFF EFPGA_CCFF_81_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_80_Q),
		.Q(EFPGA_CCFF_81_Q),
		.CFGQN(mem_outb[81]),
		.CFGQ(mem_out[81]));

	EFPGA_CCFF EFPGA_CCFF_82_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_81_Q),
		.Q(EFPGA_CCFF_82_Q),
		.CFGQN(mem_outb[82]),
		.CFGQ(mem_out[82]));

	EFPGA_CCFF EFPGA_CCFF_83_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_82_Q),
		.Q(EFPGA_CCFF_83_Q),
		.CFGQN(mem_outb[83]),
		.CFGQ(mem_out[83]));

	EFPGA_CCFF EFPGA_CCFF_84_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_83_Q),
		.Q(EFPGA_CCFF_84_Q),
		.CFGQN(mem_outb[84]),
		.CFGQ(mem_out[84]));

	EFPGA_CCFF EFPGA_CCFF_85_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_84_Q),
		.Q(EFPGA_CCFF_85_Q),
		.CFGQN(mem_outb[85]),
		.CFGQ(mem_out[85]));

	EFPGA_CCFF EFPGA_CCFF_86_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_85_Q),
		.Q(EFPGA_CCFF_86_Q),
		.CFGQN(mem_outb[86]),
		.CFGQ(mem_out[86]));

	EFPGA_CCFF EFPGA_CCFF_87_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_86_Q),
		.Q(EFPGA_CCFF_87_Q),
		.CFGQN(mem_outb[87]),
		.CFGQ(mem_out[87]));

	EFPGA_CCFF EFPGA_CCFF_88_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_87_Q),
		.Q(EFPGA_CCFF_88_Q),
		.CFGQN(mem_outb[88]),
		.CFGQ(mem_out[88]));

	EFPGA_CCFF EFPGA_CCFF_89_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_88_Q),
		.Q(EFPGA_CCFF_89_Q),
		.CFGQN(mem_outb[89]),
		.CFGQ(mem_out[89]));

	EFPGA_CCFF EFPGA_CCFF_90_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_89_Q),
		.Q(EFPGA_CCFF_90_Q),
		.CFGQN(mem_outb[90]),
		.CFGQ(mem_out[90]));

	EFPGA_CCFF EFPGA_CCFF_91_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_90_Q),
		.Q(EFPGA_CCFF_91_Q),
		.CFGQN(mem_outb[91]),
		.CFGQ(mem_out[91]));

	EFPGA_CCFF EFPGA_CCFF_92_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_91_Q),
		.Q(EFPGA_CCFF_92_Q),
		.CFGQN(mem_outb[92]),
		.CFGQ(mem_out[92]));

	EFPGA_CCFF EFPGA_CCFF_93_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_92_Q),
		.Q(EFPGA_CCFF_93_Q),
		.CFGQN(mem_outb[93]),
		.CFGQ(mem_out[93]));

	EFPGA_CCFF EFPGA_CCFF_94_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_93_Q),
		.Q(EFPGA_CCFF_94_Q),
		.CFGQN(mem_outb[94]),
		.CFGQ(mem_out[94]));

	EFPGA_CCFF EFPGA_CCFF_95_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_94_Q),
		.Q(EFPGA_CCFF_95_Q),
		.CFGQN(mem_outb[95]),
		.CFGQ(mem_out[95]));

	EFPGA_CCFF EFPGA_CCFF_96_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_95_Q),
		.Q(EFPGA_CCFF_96_Q),
		.CFGQN(mem_outb[96]),
		.CFGQ(mem_out[96]));

	EFPGA_CCFF EFPGA_CCFF_97_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_96_Q),
		.Q(EFPGA_CCFF_97_Q),
		.CFGQN(mem_outb[97]),
		.CFGQ(mem_out[97]));

	EFPGA_CCFF EFPGA_CCFF_98_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_97_Q),
		.Q(EFPGA_CCFF_98_Q),
		.CFGQN(mem_outb[98]),
		.CFGQ(mem_out[98]));

	EFPGA_CCFF EFPGA_CCFF_99_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_98_Q),
		.Q(EFPGA_CCFF_99_Q),
		.CFGQN(mem_outb[99]),
		.CFGQ(mem_out[99]));

	EFPGA_CCFF EFPGA_CCFF_100_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_99_Q),
		.Q(EFPGA_CCFF_100_Q),
		.CFGQN(mem_outb[100]),
		.CFGQ(mem_out[100]));

	EFPGA_CCFF EFPGA_CCFF_101_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_100_Q),
		.Q(EFPGA_CCFF_101_Q),
		.CFGQN(mem_outb[101]),
		.CFGQ(mem_out[101]));

	EFPGA_CCFF EFPGA_CCFF_102_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_101_Q),
		.Q(EFPGA_CCFF_102_Q),
		.CFGQN(mem_outb[102]),
		.CFGQ(mem_out[102]));

	EFPGA_CCFF EFPGA_CCFF_103_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_102_Q),
		.Q(EFPGA_CCFF_103_Q),
		.CFGQN(mem_outb[103]),
		.CFGQ(mem_out[103]));

	EFPGA_CCFF EFPGA_CCFF_104_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_103_Q),
		.Q(EFPGA_CCFF_104_Q),
		.CFGQN(mem_outb[104]),
		.CFGQ(mem_out[104]));

	EFPGA_CCFF EFPGA_CCFF_105_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_104_Q),
		.Q(EFPGA_CCFF_105_Q),
		.CFGQN(mem_outb[105]),
		.CFGQ(mem_out[105]));

	EFPGA_CCFF EFPGA_CCFF_106_ (
		.CFGE(config_enable),
		.RESET_B(prog_reset),
		.CLK(prog_clk),
		.D(EFPGA_CCFF_105_Q),
		.Q(ccff_tail),
		.CFGQN(mem_outb[106]),
		.CFGQ(mem_out[106]));

endmodule
// ----- END Verilog module for pcnt_wrapper_EFPGA_CCFF_mem -----




// ----- Verilog module for pcnt_wrapper_feedthrough_EFPGA_CCFF_mem -----
module pcnt_wrapper_feedthrough_EFPGA_CCFF_mem(feedthrough_mem_in,
                                               feedthrough_mem_inb,
                                               mem_out,
                                               mem_outb);
//----- INPUT PORTS -----
input [0:106] feedthrough_mem_in;
//----- INPUT PORTS -----
input [0:106] feedthrough_mem_inb;
//----- OUTPUT PORTS -----
output [0:106] mem_out;
//----- OUTPUT PORTS -----
output [0:106] mem_outb;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[0] = feedthrough_mem_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[1] = feedthrough_mem_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[2] = feedthrough_mem_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[3] = feedthrough_mem_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[4] = feedthrough_mem_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[5] = feedthrough_mem_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[6] = feedthrough_mem_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[7] = feedthrough_mem_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[8] = feedthrough_mem_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[9] = feedthrough_mem_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[10] = feedthrough_mem_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[11] = feedthrough_mem_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[12] = feedthrough_mem_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[13] = feedthrough_mem_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[14] = feedthrough_mem_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[15] = feedthrough_mem_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[16] = feedthrough_mem_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[17] = feedthrough_mem_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[18] = feedthrough_mem_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[19] = feedthrough_mem_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[20] = feedthrough_mem_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[21] = feedthrough_mem_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[22] = feedthrough_mem_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[23] = feedthrough_mem_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[24] = feedthrough_mem_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[25] = feedthrough_mem_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[26] = feedthrough_mem_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[27] = feedthrough_mem_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[28] = feedthrough_mem_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[29] = feedthrough_mem_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[30] = feedthrough_mem_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[31] = feedthrough_mem_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[32] = feedthrough_mem_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[33] = feedthrough_mem_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[34] = feedthrough_mem_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[35] = feedthrough_mem_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[36] = feedthrough_mem_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[37] = feedthrough_mem_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[38] = feedthrough_mem_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[39] = feedthrough_mem_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[40] = feedthrough_mem_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[41] = feedthrough_mem_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[42] = feedthrough_mem_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[43] = feedthrough_mem_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[44] = feedthrough_mem_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[45] = feedthrough_mem_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[46] = feedthrough_mem_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[47] = feedthrough_mem_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[48] = feedthrough_mem_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[49] = feedthrough_mem_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[50] = feedthrough_mem_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[51] = feedthrough_mem_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[52] = feedthrough_mem_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[53] = feedthrough_mem_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[54] = feedthrough_mem_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[55] = feedthrough_mem_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[56] = feedthrough_mem_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[57] = feedthrough_mem_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[58] = feedthrough_mem_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[59] = feedthrough_mem_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[60] = feedthrough_mem_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[61] = feedthrough_mem_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[62] = feedthrough_mem_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[63] = feedthrough_mem_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[64] = feedthrough_mem_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[65] = feedthrough_mem_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[66] = feedthrough_mem_in[66];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[67] = feedthrough_mem_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[68] = feedthrough_mem_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[69] = feedthrough_mem_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[70] = feedthrough_mem_in[70];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[71] = feedthrough_mem_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[72] = feedthrough_mem_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[73] = feedthrough_mem_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[74] = feedthrough_mem_in[74];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[75] = feedthrough_mem_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[76] = feedthrough_mem_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[77] = feedthrough_mem_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[78] = feedthrough_mem_in[78];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[79] = feedthrough_mem_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[80] = feedthrough_mem_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[81] = feedthrough_mem_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[82] = feedthrough_mem_in[82];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[83] = feedthrough_mem_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[84] = feedthrough_mem_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[85] = feedthrough_mem_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[86] = feedthrough_mem_in[86];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[87] = feedthrough_mem_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[88] = feedthrough_mem_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[89] = feedthrough_mem_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[90] = feedthrough_mem_in[90];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[91] = feedthrough_mem_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[92] = feedthrough_mem_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[93] = feedthrough_mem_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[94] = feedthrough_mem_in[94];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[95] = feedthrough_mem_in[95];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[96] = feedthrough_mem_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[97] = feedthrough_mem_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[98] = feedthrough_mem_in[98];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[99] = feedthrough_mem_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[100] = feedthrough_mem_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[101] = feedthrough_mem_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[102] = feedthrough_mem_in[102];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[103] = feedthrough_mem_in[103];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[104] = feedthrough_mem_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[105] = feedthrough_mem_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_out[106] = feedthrough_mem_in[106];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[0] = feedthrough_mem_inb[0];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[1] = feedthrough_mem_inb[1];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[2] = feedthrough_mem_inb[2];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[3] = feedthrough_mem_inb[3];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[4] = feedthrough_mem_inb[4];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[5] = feedthrough_mem_inb[5];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[6] = feedthrough_mem_inb[6];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[7] = feedthrough_mem_inb[7];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[8] = feedthrough_mem_inb[8];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[9] = feedthrough_mem_inb[9];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[10] = feedthrough_mem_inb[10];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[11] = feedthrough_mem_inb[11];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[12] = feedthrough_mem_inb[12];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[13] = feedthrough_mem_inb[13];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[14] = feedthrough_mem_inb[14];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[15] = feedthrough_mem_inb[15];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[16] = feedthrough_mem_inb[16];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[17] = feedthrough_mem_inb[17];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[18] = feedthrough_mem_inb[18];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[19] = feedthrough_mem_inb[19];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[20] = feedthrough_mem_inb[20];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[21] = feedthrough_mem_inb[21];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[22] = feedthrough_mem_inb[22];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[23] = feedthrough_mem_inb[23];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[24] = feedthrough_mem_inb[24];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[25] = feedthrough_mem_inb[25];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[26] = feedthrough_mem_inb[26];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[27] = feedthrough_mem_inb[27];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[28] = feedthrough_mem_inb[28];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[29] = feedthrough_mem_inb[29];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[30] = feedthrough_mem_inb[30];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[31] = feedthrough_mem_inb[31];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[32] = feedthrough_mem_inb[32];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[33] = feedthrough_mem_inb[33];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[34] = feedthrough_mem_inb[34];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[35] = feedthrough_mem_inb[35];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[36] = feedthrough_mem_inb[36];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[37] = feedthrough_mem_inb[37];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[38] = feedthrough_mem_inb[38];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[39] = feedthrough_mem_inb[39];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[40] = feedthrough_mem_inb[40];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[41] = feedthrough_mem_inb[41];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[42] = feedthrough_mem_inb[42];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[43] = feedthrough_mem_inb[43];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[44] = feedthrough_mem_inb[44];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[45] = feedthrough_mem_inb[45];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[46] = feedthrough_mem_inb[46];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[47] = feedthrough_mem_inb[47];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[48] = feedthrough_mem_inb[48];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[49] = feedthrough_mem_inb[49];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[50] = feedthrough_mem_inb[50];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[51] = feedthrough_mem_inb[51];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[52] = feedthrough_mem_inb[52];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[53] = feedthrough_mem_inb[53];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[54] = feedthrough_mem_inb[54];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[55] = feedthrough_mem_inb[55];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[56] = feedthrough_mem_inb[56];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[57] = feedthrough_mem_inb[57];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[58] = feedthrough_mem_inb[58];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[59] = feedthrough_mem_inb[59];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[60] = feedthrough_mem_inb[60];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[61] = feedthrough_mem_inb[61];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[62] = feedthrough_mem_inb[62];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[63] = feedthrough_mem_inb[63];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[64] = feedthrough_mem_inb[64];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[65] = feedthrough_mem_inb[65];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[66] = feedthrough_mem_inb[66];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[67] = feedthrough_mem_inb[67];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[68] = feedthrough_mem_inb[68];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[69] = feedthrough_mem_inb[69];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[70] = feedthrough_mem_inb[70];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[71] = feedthrough_mem_inb[71];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[72] = feedthrough_mem_inb[72];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[73] = feedthrough_mem_inb[73];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[74] = feedthrough_mem_inb[74];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[75] = feedthrough_mem_inb[75];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[76] = feedthrough_mem_inb[76];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[77] = feedthrough_mem_inb[77];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[78] = feedthrough_mem_inb[78];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[79] = feedthrough_mem_inb[79];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[80] = feedthrough_mem_inb[80];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[81] = feedthrough_mem_inb[81];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[82] = feedthrough_mem_inb[82];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[83] = feedthrough_mem_inb[83];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[84] = feedthrough_mem_inb[84];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[85] = feedthrough_mem_inb[85];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[86] = feedthrough_mem_inb[86];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[87] = feedthrough_mem_inb[87];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[88] = feedthrough_mem_inb[88];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[89] = feedthrough_mem_inb[89];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[90] = feedthrough_mem_inb[90];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[91] = feedthrough_mem_inb[91];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[92] = feedthrough_mem_inb[92];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[93] = feedthrough_mem_inb[93];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[94] = feedthrough_mem_inb[94];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[95] = feedthrough_mem_inb[95];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[96] = feedthrough_mem_inb[96];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[97] = feedthrough_mem_inb[97];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[98] = feedthrough_mem_inb[98];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[99] = feedthrough_mem_inb[99];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[100] = feedthrough_mem_inb[100];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[101] = feedthrough_mem_inb[101];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[102] = feedthrough_mem_inb[102];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[103] = feedthrough_mem_inb[103];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[104] = feedthrough_mem_inb[104];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[105] = feedthrough_mem_inb[105];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign mem_outb[106] = feedthrough_mem_inb[106];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

endmodule
// ----- END Verilog module for pcnt_wrapper_feedthrough_EFPGA_CCFF_mem -----




// ----- Verilog module for grid_clb_config_group_mem_size885 -----
module grid_clb_config_group_mem_size885(config_enable,
                                         prog_reset,
                                         prog_clk,
                                         ccff_head,
                                         mem_out,
                                         mem_outb,
                                         ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:884] mem_out;
//----- OUTPUT PORTS -----
output [0:884] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[0:32]),
		.mem_outb(mem_outb[0:32]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_0_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[47:79]),
		.mem_outb(mem_outb[47:79]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_1_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[94:126]),
		.mem_outb(mem_outb[94:126]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_2_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[141:173]),
		.mem_outb(mem_outb[141:173]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_3_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[188:220]),
		.mem_outb(mem_outb[188:220]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_4_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[235:267]),
		.mem_outb(mem_outb[235:267]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_5_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[282:314]),
		.mem_outb(mem_outb[282:314]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_6_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[329:361]),
		.mem_outb(mem_outb[329:361]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_8_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_7_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_8_ccff_tail),
		.mem_out(mem_out[376:408]),
		.mem_outb(mem_outb[376:408]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_9_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_8_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_9_ccff_tail),
		.mem_out(mem_out[423:455]),
		.mem_outb(mem_outb[423:455]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_10_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_9_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_10_ccff_tail),
		.mem_out(mem_out[470:502]),
		.mem_outb(mem_outb[470:502]));

	frac_lut5_arith_EFPGA_CCFF_mem frac_lut5_arith_EFPGA_CCFF_mem_11_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_10_ccff_tail),
		.ccff_tail(frac_lut5_arith_EFPGA_CCFF_mem_11_ccff_tail),
		.mem_out(mem_out[517:549]),
		.mem_outb(mem_outb[517:549]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_0_ccff_tail),
		.mem_out(mem_out[33]),
		.mem_outb(mem_outb[33]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_1_ccff_tail),
		.mem_out(mem_out[80]),
		.mem_outb(mem_outb[80]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_2_ccff_tail),
		.mem_out(mem_out[127]),
		.mem_outb(mem_outb[127]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_3_ccff_tail),
		.mem_out(mem_out[174]),
		.mem_outb(mem_outb[174]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_4_ccff_tail),
		.mem_out(mem_out[221]),
		.mem_outb(mem_outb[221]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_5_ccff_tail),
		.mem_out(mem_out[268]),
		.mem_outb(mem_outb[268]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_6_ccff_tail),
		.mem_out(mem_out[315]),
		.mem_outb(mem_outb[315]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_7_ccff_tail),
		.mem_out(mem_out[362]),
		.mem_outb(mem_outb[362]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_8_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_8_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_8_ccff_tail),
		.mem_out(mem_out[409]),
		.mem_outb(mem_outb[409]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_9_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_9_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_9_ccff_tail),
		.mem_out(mem_out[456]),
		.mem_outb(mem_outb[456]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_10_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_10_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_10_ccff_tail),
		.mem_out(mem_out[503]),
		.mem_outb(mem_outb[503]));

	pb_mux_no_const_input_size2_mem mem_frac_logic_out_0_11_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(frac_lut5_arith_EFPGA_CCFF_mem_11_ccff_tail),
		.ccff_tail(pb_mux_no_const_input_size2_mem_11_ccff_tail),
		.mem_out(mem_out[550]),
		.mem_outb(mem_outb[550]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_0_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[34:37]),
		.mem_outb(mem_outb[34:37]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[38:41]),
		.mem_outb(mem_outb[38:41]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_1_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[81:84]),
		.mem_outb(mem_outb[81:84]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[85:88]),
		.mem_outb(mem_outb[85:88]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_2_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[128:131]),
		.mem_outb(mem_outb[128:131]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[132:135]),
		.mem_outb(mem_outb[132:135]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_3_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[175:178]),
		.mem_outb(mem_outb[175:178]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[179:182]),
		.mem_outb(mem_outb[179:182]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_8_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_4_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_8_ccff_tail),
		.mem_out(mem_out[222:225]),
		.mem_outb(mem_outb[222:225]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_9_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_8_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_9_ccff_tail),
		.mem_out(mem_out[226:229]),
		.mem_outb(mem_outb[226:229]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_10_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_5_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_10_ccff_tail),
		.mem_out(mem_out[269:272]),
		.mem_outb(mem_outb[269:272]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_11_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_10_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_11_ccff_tail),
		.mem_out(mem_out[273:276]),
		.mem_outb(mem_outb[273:276]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_12_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_6_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_12_ccff_tail),
		.mem_out(mem_out[316:319]),
		.mem_outb(mem_outb[316:319]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_13_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_12_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_13_ccff_tail),
		.mem_out(mem_out[320:323]),
		.mem_outb(mem_outb[320:323]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_14_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_7_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_14_ccff_tail),
		.mem_out(mem_out[363:366]),
		.mem_outb(mem_outb[363:366]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_15_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_14_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_15_ccff_tail),
		.mem_out(mem_out[367:370]),
		.mem_outb(mem_outb[367:370]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_16_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_8_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_16_ccff_tail),
		.mem_out(mem_out[410:413]),
		.mem_outb(mem_outb[410:413]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_17_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_16_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_17_ccff_tail),
		.mem_out(mem_out[414:417]),
		.mem_outb(mem_outb[414:417]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_18_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_9_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_18_ccff_tail),
		.mem_out(mem_out[457:460]),
		.mem_outb(mem_outb[457:460]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_19_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_18_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_19_ccff_tail),
		.mem_out(mem_out[461:464]),
		.mem_outb(mem_outb[461:464]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_20_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_10_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_20_ccff_tail),
		.mem_out(mem_out[504:507]),
		.mem_outb(mem_outb[504:507]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_21_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_20_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_21_ccff_tail),
		.mem_out(mem_out[508:511]),
		.mem_outb(mem_outb[508:511]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_22_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_no_const_input_size2_mem_11_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_22_ccff_tail),
		.mem_out(mem_out[551:554]),
		.mem_outb(mem_outb[551:554]));

	mmff_wrapper_EFPGA_CCFF_mem mmff_wrapper_EFPGA_CCFF_mem_23_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_22_ccff_tail),
		.ccff_tail(mmff_wrapper_EFPGA_CCFF_mem_23_ccff_tail),
		.mem_out(mem_out[555:558]),
		.mem_outb(mem_outb[555:558]));

	pb_mux_highload_size2_mem mem_fabric_out_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_0_ccff_tail),
		.mem_out(mem_out[42]),
		.mem_outb(mem_outb[42]));

	pb_mux_highload_size2_mem mem_fabric_out_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_1_ccff_tail),
		.mem_out(mem_out[89]),
		.mem_outb(mem_outb[89]));

	pb_mux_highload_size2_mem mem_fabric_out_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_2_ccff_tail),
		.mem_out(mem_out[136]),
		.mem_outb(mem_outb[136]));

	pb_mux_highload_size2_mem mem_fabric_out_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_3_ccff_tail),
		.mem_out(mem_out[183]),
		.mem_outb(mem_outb[183]));

	pb_mux_highload_size2_mem mem_fabric_out_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_9_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_4_ccff_tail),
		.mem_out(mem_out[230]),
		.mem_outb(mem_outb[230]));

	pb_mux_highload_size2_mem mem_fabric_out_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_11_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_5_ccff_tail),
		.mem_out(mem_out[277]),
		.mem_outb(mem_outb[277]));

	pb_mux_highload_size2_mem mem_fabric_out_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_13_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_6_ccff_tail),
		.mem_out(mem_out[324]),
		.mem_outb(mem_outb[324]));

	pb_mux_highload_size2_mem mem_fabric_out_0_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_15_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_7_ccff_tail),
		.mem_out(mem_out[371]),
		.mem_outb(mem_outb[371]));

	pb_mux_highload_size2_mem mem_fabric_out_0_8_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_17_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_8_ccff_tail),
		.mem_out(mem_out[418]),
		.mem_outb(mem_outb[418]));

	pb_mux_highload_size2_mem mem_fabric_out_0_9_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_19_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_9_ccff_tail),
		.mem_out(mem_out[465]),
		.mem_outb(mem_outb[465]));

	pb_mux_highload_size2_mem mem_fabric_out_0_10_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_21_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_10_ccff_tail),
		.mem_out(mem_out[512]),
		.mem_outb(mem_outb[512]));

	pb_mux_highload_size2_mem mem_fabric_out_0_11_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmff_wrapper_EFPGA_CCFF_mem_23_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_11_ccff_tail),
		.mem_out(mem_out[559]),
		.mem_outb(mem_outb[559]));

	pb_mux_highload_size3_mem mem_fabric_out_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_0_ccff_tail),
		.mem_out(mem_out[43:44]),
		.mem_outb(mem_outb[43:44]));

	pb_mux_highload_size3_mem mem_fabric_out_1_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_1_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	pb_mux_highload_size3_mem mem_fabric_out_1_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_2_ccff_tail),
		.mem_out(mem_out[137:138]),
		.mem_outb(mem_outb[137:138]));

	pb_mux_highload_size3_mem mem_fabric_out_1_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_3_ccff_tail),
		.mem_out(mem_out[184:185]),
		.mem_outb(mem_outb[184:185]));

	pb_mux_highload_size3_mem mem_fabric_out_1_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_4_ccff_tail),
		.mem_out(mem_out[231:232]),
		.mem_outb(mem_outb[231:232]));

	pb_mux_highload_size3_mem mem_fabric_out_1_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_5_ccff_tail),
		.mem_out(mem_out[278:279]),
		.mem_outb(mem_outb[278:279]));

	pb_mux_highload_size3_mem mem_fabric_out_1_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_6_ccff_tail),
		.mem_out(mem_out[325:326]),
		.mem_outb(mem_outb[325:326]));

	pb_mux_highload_size3_mem mem_fabric_out_1_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_7_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_7_ccff_tail),
		.mem_out(mem_out[372:373]),
		.mem_outb(mem_outb[372:373]));

	pb_mux_highload_size3_mem mem_fabric_out_1_8_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_8_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_8_ccff_tail),
		.mem_out(mem_out[419:420]),
		.mem_outb(mem_outb[419:420]));

	pb_mux_highload_size3_mem mem_fabric_out_1_9_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_9_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_9_ccff_tail),
		.mem_out(mem_out[466:467]),
		.mem_outb(mem_outb[466:467]));

	pb_mux_highload_size3_mem mem_fabric_out_1_10_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_10_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_10_ccff_tail),
		.mem_out(mem_out[513:514]),
		.mem_outb(mem_outb[513:514]));

	pb_mux_highload_size3_mem mem_fabric_out_1_11_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_11_ccff_tail),
		.ccff_tail(pb_mux_highload_size3_mem_11_ccff_tail),
		.mem_out(mem_out[560:561]),
		.mem_outb(mem_outb[560:561]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_0_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_0_ccff_tail),
		.mem_out(mem_out[45:46]),
		.mem_outb(mem_outb[45:46]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_1_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_1_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_2_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_2_ccff_tail),
		.mem_out(mem_out[139:140]),
		.mem_outb(mem_outb[139:140]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_3_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_3_ccff_tail),
		.mem_out(mem_out[186:187]),
		.mem_outb(mem_outb[186:187]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_4_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_4_ccff_tail),
		.mem_out(mem_out[233:234]),
		.mem_outb(mem_outb[233:234]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_5_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_5_ccff_tail),
		.mem_out(mem_out[280:281]),
		.mem_outb(mem_outb[280:281]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_6_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_6_ccff_tail),
		.mem_out(mem_out[327:328]),
		.mem_outb(mem_outb[327:328]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_7_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_7_ccff_tail),
		.mem_out(mem_out[374:375]),
		.mem_outb(mem_outb[374:375]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_8_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_8_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_8_ccff_tail),
		.mem_out(mem_out[421:422]),
		.mem_outb(mem_outb[421:422]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_9_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_9_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_9_ccff_tail),
		.mem_out(mem_out[468:469]),
		.mem_outb(mem_outb[468:469]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_10_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_10_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_10_ccff_tail),
		.mem_out(mem_out[515:516]),
		.mem_outb(mem_outb[515:516]));

	pb_mux_size2_mem mem_p_ff_p_ff_1_D_0_11_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size3_mem_11_ccff_tail),
		.ccff_tail(pb_mux_size2_mem_11_ccff_tail),
		.mem_out(mem_out[562:563]),
		.mem_outb(mem_outb[562:563]));

	pcnt_wrapper_EFPGA_CCFF_mem pcnt_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_size2_mem_11_ccff_tail),
		.ccff_tail(pcnt_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[564:670]),
		.mem_outb(mem_outb[564:670]));

	pcnt_wrapper_EFPGA_CCFF_mem pcnt_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pcnt_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pcnt_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[671:777]),
		.mem_outb(mem_outb[671:777]));

	pcnt_wrapper_EFPGA_CCFF_mem pcnt_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pcnt_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[778:884]),
		.mem_outb(mem_outb[778:884]));

endmodule
// ----- END Verilog module for grid_clb_config_group_mem_size885 -----




// ----- Verilog module for grid_io_bottomL_bottom_config_group_mem_size140 -----
module grid_io_bottomL_bottom_config_group_mem_size140(config_enable,
                                                       prog_reset,
                                                       prog_clk,
                                                       ccff_head,
                                                       mem_out,
                                                       mem_outb,
                                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:139] mem_out;
//----- OUTPUT PORTS -----
output [0:139] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	pinput_dchain_extmode_EFPGA_CCFF_mem pinput_dchain_extmode_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(pinput_dchain_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[0:4]),
		.mem_outb(mem_outb[0:4]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_dchain_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[5:11]),
		.mem_outb(mem_outb[5:11]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[14:20]),
		.mem_outb(mem_outb[14:20]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[23:29]),
		.mem_outb(mem_outb[23:29]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[32:38]),
		.mem_outb(mem_outb[32:38]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[41:47]),
		.mem_outb(mem_outb[41:47]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[50:56]),
		.mem_outb(mem_outb[50:56]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[59:65]),
		.mem_outb(mem_outb[59:65]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[68:74]),
		.mem_outb(mem_outb[68:74]));

	pb_mux_highload_size2_mem mem_pi_pdc_ecb1_pad_a2f_o_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_0_ccff_tail),
		.mem_out(mem_out[12]),
		.mem_outb(mem_outb[12]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_1_ccff_tail),
		.mem_out(mem_out[21]),
		.mem_outb(mem_outb[21]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_2_ccff_tail),
		.mem_out(mem_out[30]),
		.mem_outb(mem_outb[30]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_3_ccff_tail),
		.mem_out(mem_out[39]),
		.mem_outb(mem_outb[39]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_4_ccff_tail),
		.mem_out(mem_out[48]),
		.mem_outb(mem_outb[48]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_5_ccff_tail),
		.mem_out(mem_out[57]),
		.mem_outb(mem_outb[57]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_6_ccff_tail),
		.mem_out(mem_out[66]),
		.mem_outb(mem_outb[66]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_7_ccff_tail),
		.mem_out(mem_out[75]),
		.mem_outb(mem_outb[75]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_8_ccff_tail),
		.mem_out(mem_out[83]),
		.mem_outb(mem_outb[83]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_9_ccff_tail),
		.mem_out(mem_out[91]),
		.mem_outb(mem_outb[91]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_10_ccff_tail),
		.mem_out(mem_out[99]),
		.mem_outb(mem_outb[99]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_11_ccff_tail),
		.mem_out(mem_out[107]),
		.mem_outb(mem_outb[107]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_12_ccff_tail),
		.mem_out(mem_out[115]),
		.mem_outb(mem_outb[115]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_13_ccff_tail),
		.mem_out(mem_out[123]),
		.mem_outb(mem_outb[123]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_14_ccff_tail),
		.mem_out(mem_out[131]),
		.mem_outb(mem_outb[131]));

	pb_mux_highload_size2_mem mem_io_po_cko_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[139]),
		.mem_outb(mem_outb[139]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_0_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[13]),
		.mem_outb(mem_outb[13]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_1_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[22]),
		.mem_outb(mem_outb[22]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_2_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[31]),
		.mem_outb(mem_outb[31]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_3_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[40]),
		.mem_outb(mem_outb[40]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_4_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[49]),
		.mem_outb(mem_outb[49]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_5_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[58]),
		.mem_outb(mem_outb[58]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_6_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[67]),
		.mem_outb(mem_outb[67]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_7_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[76:82]),
		.mem_outb(mem_outb[76:82]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_8_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[84:90]),
		.mem_outb(mem_outb[84:90]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_9_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[92:98]),
		.mem_outb(mem_outb[92:98]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_10_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[100:106]),
		.mem_outb(mem_outb[100:106]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_11_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[108:114]),
		.mem_outb(mem_outb[108:114]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_12_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[116:122]),
		.mem_outb(mem_outb[116:122]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_13_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[124:130]),
		.mem_outb(mem_outb[124:130]));

	mmffosc2cko_wrapper_EFPGA_CCFF_mem mmffosc2cko_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_14_ccff_tail),
		.ccff_tail(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[132:138]),
		.mem_outb(mem_outb[132:138]));

endmodule
// ----- END Verilog module for grid_io_bottomL_bottom_config_group_mem_size140 -----




// ----- Verilog module for grid_io_leftL_left_config_group_mem_size136 -----
module grid_io_leftL_left_config_group_mem_size136(config_enable,
                                                   prog_reset,
                                                   prog_clk,
                                                   ccff_head,
                                                   mem_out,
                                                   mem_outb,
                                                   ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:135] mem_out;
//----- OUTPUT PORTS -----
output [0:135] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[0]),
		.mem_outb(mem_outb[0]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_0_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[9]),
		.mem_outb(mem_outb[9]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_1_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[18]),
		.mem_outb(mem_outb[18]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_2_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[27]),
		.mem_outb(mem_outb[27]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_3_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[36]),
		.mem_outb(mem_outb[36]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_4_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[45]),
		.mem_outb(mem_outb[45]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_5_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[54]),
		.mem_outb(mem_outb[54]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_6_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[63]),
		.mem_outb(mem_outb[63]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[1:7]),
		.mem_outb(mem_outb[1:7]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[10:16]),
		.mem_outb(mem_outb[10:16]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[19:25]),
		.mem_outb(mem_outb[19:25]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[28:34]),
		.mem_outb(mem_outb[28:34]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[37:43]),
		.mem_outb(mem_outb[37:43]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[46:52]),
		.mem_outb(mem_outb[46:52]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[55:61]),
		.mem_outb(mem_outb[55:61]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[64:70]),
		.mem_outb(mem_outb[64:70]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_0_ccff_tail),
		.mem_out(mem_out[8]),
		.mem_outb(mem_outb[8]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_1_ccff_tail),
		.mem_out(mem_out[17]),
		.mem_outb(mem_outb[17]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_2_ccff_tail),
		.mem_out(mem_out[26]),
		.mem_outb(mem_outb[26]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_3_ccff_tail),
		.mem_out(mem_out[35]),
		.mem_outb(mem_outb[35]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_4_ccff_tail),
		.mem_out(mem_out[44]),
		.mem_outb(mem_outb[44]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_5_ccff_tail),
		.mem_out(mem_out[53]),
		.mem_outb(mem_outb[53]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_6_ccff_tail),
		.mem_out(mem_out[62]),
		.mem_outb(mem_outb[62]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_7_ccff_tail),
		.mem_out(mem_out[71]),
		.mem_outb(mem_outb[71]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_8_ccff_tail),
		.mem_out(mem_out[79]),
		.mem_outb(mem_outb[79]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_9_ccff_tail),
		.mem_out(mem_out[87]),
		.mem_outb(mem_outb[87]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_10_ccff_tail),
		.mem_out(mem_out[95]),
		.mem_outb(mem_outb[95]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_11_ccff_tail),
		.mem_out(mem_out[103]),
		.mem_outb(mem_outb[103]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_12_ccff_tail),
		.mem_out(mem_out[111]),
		.mem_outb(mem_outb[111]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_13_ccff_tail),
		.mem_out(mem_out[119]),
		.mem_outb(mem_outb[119]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_14_ccff_tail),
		.mem_out(mem_out[127]),
		.mem_outb(mem_outb[127]));

	pb_mux_highload_size2_mem mem_io_po_cko_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[135]),
		.mem_outb(mem_outb[135]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_7_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[72:78]),
		.mem_outb(mem_outb[72:78]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_8_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[80:86]),
		.mem_outb(mem_outb[80:86]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_9_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[88:94]),
		.mem_outb(mem_outb[88:94]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_10_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[96:102]),
		.mem_outb(mem_outb[96:102]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_11_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[104:110]),
		.mem_outb(mem_outb[104:110]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_12_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[112:118]),
		.mem_outb(mem_outb[112:118]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_13_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[120:126]),
		.mem_outb(mem_outb[120:126]));

	mmffosc2cko_wrapper_EFPGA_CCFF_mem mmffosc2cko_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_14_ccff_tail),
		.ccff_tail(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[128:134]),
		.mem_outb(mem_outb[128:134]));

endmodule
// ----- END Verilog module for grid_io_leftL_left_config_group_mem_size136 -----




// ----- Verilog module for grid_io_rightL_right_config_group_mem_size136 -----
module grid_io_rightL_right_config_group_mem_size136(config_enable,
                                                     prog_reset,
                                                     prog_clk,
                                                     ccff_head,
                                                     mem_out,
                                                     mem_outb,
                                                     ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:135] mem_out;
//----- OUTPUT PORTS -----
output [0:135] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[0]),
		.mem_outb(mem_outb[0]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_0_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[9]),
		.mem_outb(mem_outb[9]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_1_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[18]),
		.mem_outb(mem_outb[18]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_2_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[27]),
		.mem_outb(mem_outb[27]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_3_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[36]),
		.mem_outb(mem_outb[36]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_4_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[45]),
		.mem_outb(mem_outb[45]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_5_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[54]),
		.mem_outb(mem_outb[54]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_6_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[63]),
		.mem_outb(mem_outb[63]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[1:7]),
		.mem_outb(mem_outb[1:7]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[10:16]),
		.mem_outb(mem_outb[10:16]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[19:25]),
		.mem_outb(mem_outb[19:25]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[28:34]),
		.mem_outb(mem_outb[28:34]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[37:43]),
		.mem_outb(mem_outb[37:43]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[46:52]),
		.mem_outb(mem_outb[46:52]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[55:61]),
		.mem_outb(mem_outb[55:61]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[64:70]),
		.mem_outb(mem_outb[64:70]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_0_ccff_tail),
		.mem_out(mem_out[8]),
		.mem_outb(mem_outb[8]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_1_ccff_tail),
		.mem_out(mem_out[17]),
		.mem_outb(mem_outb[17]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_2_ccff_tail),
		.mem_out(mem_out[26]),
		.mem_outb(mem_outb[26]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_3_ccff_tail),
		.mem_out(mem_out[35]),
		.mem_outb(mem_outb[35]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_4_ccff_tail),
		.mem_out(mem_out[44]),
		.mem_outb(mem_outb[44]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_5_ccff_tail),
		.mem_out(mem_out[53]),
		.mem_outb(mem_outb[53]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_6_ccff_tail),
		.mem_out(mem_out[62]),
		.mem_outb(mem_outb[62]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_7_ccff_tail),
		.mem_out(mem_out[71]),
		.mem_outb(mem_outb[71]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_8_ccff_tail),
		.mem_out(mem_out[79]),
		.mem_outb(mem_outb[79]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_9_ccff_tail),
		.mem_out(mem_out[87]),
		.mem_outb(mem_outb[87]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_10_ccff_tail),
		.mem_out(mem_out[95]),
		.mem_outb(mem_outb[95]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_11_ccff_tail),
		.mem_out(mem_out[103]),
		.mem_outb(mem_outb[103]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_12_ccff_tail),
		.mem_out(mem_out[111]),
		.mem_outb(mem_outb[111]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_13_ccff_tail),
		.mem_out(mem_out[119]),
		.mem_outb(mem_outb[119]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_14_ccff_tail),
		.mem_out(mem_out[127]),
		.mem_outb(mem_outb[127]));

	pb_mux_highload_size2_mem mem_io_po_cko_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[135]),
		.mem_outb(mem_outb[135]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_7_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[72:78]),
		.mem_outb(mem_outb[72:78]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_8_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[80:86]),
		.mem_outb(mem_outb[80:86]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_9_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[88:94]),
		.mem_outb(mem_outb[88:94]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_10_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[96:102]),
		.mem_outb(mem_outb[96:102]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_11_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[104:110]),
		.mem_outb(mem_outb[104:110]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_12_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[112:118]),
		.mem_outb(mem_outb[112:118]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_13_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[120:126]),
		.mem_outb(mem_outb[120:126]));

	mmffosc2cko_wrapper_EFPGA_CCFF_mem mmffosc2cko_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_14_ccff_tail),
		.ccff_tail(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[128:134]),
		.mem_outb(mem_outb[128:134]));

endmodule
// ----- END Verilog module for grid_io_rightL_right_config_group_mem_size136 -----




// ----- Verilog module for grid_io_topL_top_config_group_mem_size136 -----
module grid_io_topL_top_config_group_mem_size136(config_enable,
                                                 prog_reset,
                                                 prog_clk,
                                                 ccff_head,
                                                 mem_out,
                                                 mem_outb,
                                                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:135] mem_out;
//----- OUTPUT PORTS -----
output [0:135] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[0]),
		.mem_outb(mem_outb[0]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_0_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[9]),
		.mem_outb(mem_outb[9]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_1_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[18]),
		.mem_outb(mem_outb[18]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_2_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[27]),
		.mem_outb(mem_outb[27]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_3_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[36]),
		.mem_outb(mem_outb[36]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_4_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[45]),
		.mem_outb(mem_outb[45]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_5_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[54]),
		.mem_outb(mem_outb[54]));

	pinput_extmode_EFPGA_CCFF_mem pinput_extmode_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_6_ccff_tail),
		.ccff_tail(pinput_extmode_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[63]),
		.mem_outb(mem_outb[63]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[1:7]),
		.mem_outb(mem_outb[1:7]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[10:16]),
		.mem_outb(mem_outb[10:16]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[19:25]),
		.mem_outb(mem_outb[19:25]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[28:34]),
		.mem_outb(mem_outb[28:34]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[37:43]),
		.mem_outb(mem_outb[37:43]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[46:52]),
		.mem_outb(mem_outb[46:52]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[55:61]),
		.mem_outb(mem_outb[55:61]));

	mmffisc2_wrapper_EFPGA_CCFF_mem mmffisc2_wrapper_EFPGA_CCFF_mem_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pinput_extmode_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.mem_out(mem_out[64:70]),
		.mem_outb(mem_outb[64:70]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_0_ccff_tail),
		.mem_out(mem_out[8]),
		.mem_outb(mem_outb[8]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_1_ccff_tail),
		.mem_out(mem_out[17]),
		.mem_outb(mem_outb[17]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_2_ccff_tail),
		.mem_out(mem_out[26]),
		.mem_outb(mem_outb[26]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_3_ccff_tail),
		.mem_out(mem_out[35]),
		.mem_outb(mem_outb[35]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_4_ccff_tail),
		.mem_out(mem_out[44]),
		.mem_outb(mem_outb[44]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_5_ccff_tail),
		.mem_out(mem_out[53]),
		.mem_outb(mem_outb[53]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_6_ccff_tail),
		.mem_out(mem_out[62]),
		.mem_outb(mem_outb[62]));

	pb_mux_highload_size2_mem mem_pi_pad_a2f_o_0_7_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffisc2_wrapper_EFPGA_CCFF_mem_7_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_7_ccff_tail),
		.mem_out(mem_out[71]),
		.mem_outb(mem_outb[71]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_8_ccff_tail),
		.mem_out(mem_out[79]),
		.mem_outb(mem_outb[79]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_9_ccff_tail),
		.mem_out(mem_out[87]),
		.mem_outb(mem_outb[87]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_10_ccff_tail),
		.mem_out(mem_out[95]),
		.mem_outb(mem_outb[95]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_11_ccff_tail),
		.mem_out(mem_out[103]),
		.mem_outb(mem_outb[103]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_12_ccff_tail),
		.mem_out(mem_out[111]),
		.mem_outb(mem_outb[111]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_13_ccff_tail),
		.mem_out(mem_out[119]),
		.mem_outb(mem_outb[119]));

	pb_mux_highload_size2_mem mem_io_po_core_0_outpad_0_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.ccff_tail(pb_mux_highload_size2_mem_14_ccff_tail),
		.mem_out(mem_out[127]),
		.mem_outb(mem_outb[127]));

	pb_mux_highload_size2_mem mem_io_po_cko_core_0_outpad_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[135]),
		.mem_outb(mem_outb[135]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_7_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[72:78]),
		.mem_outb(mem_outb[72:78]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_1_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_8_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_1_ccff_tail),
		.mem_out(mem_out[80:86]),
		.mem_outb(mem_outb[80:86]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_2_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_9_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_2_ccff_tail),
		.mem_out(mem_out[88:94]),
		.mem_outb(mem_outb[88:94]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_3_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_10_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_3_ccff_tail),
		.mem_out(mem_out[96:102]),
		.mem_outb(mem_outb[96:102]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_4_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_11_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_4_ccff_tail),
		.mem_out(mem_out[104:110]),
		.mem_outb(mem_outb[104:110]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_5_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_12_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_5_ccff_tail),
		.mem_out(mem_out[112:118]),
		.mem_outb(mem_outb[112:118]));

	mmffosc2_wrapper_EFPGA_CCFF_mem mmffosc2_wrapper_EFPGA_CCFF_mem_6_ (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_13_ccff_tail),
		.ccff_tail(mmffosc2_wrapper_EFPGA_CCFF_mem_6_ccff_tail),
		.mem_out(mem_out[120:126]),
		.mem_outb(mem_outb[120:126]));

	mmffosc2cko_wrapper_EFPGA_CCFF_mem mmffosc2cko_wrapper_EFPGA_CCFF_mem (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(pb_mux_highload_size2_mem_14_ccff_tail),
		.ccff_tail(mmffosc2cko_wrapper_EFPGA_CCFF_mem_0_ccff_tail),
		.mem_out(mem_out[128:134]),
		.mem_outb(mem_outb[128:134]));

endmodule
// ----- END Verilog module for grid_io_topL_top_config_group_mem_size136 -----




// ----- Verilog module for sb_0__config_group_mem_size265 -----
module sb_0__config_group_mem_size265(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:264] mem_out;
//----- OUTPUT PORTS -----
output [0:264] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size6_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size6_mem_0_ccff_tail),
		.mem_out(mem_out[0:2]),
		.mem_outb(mem_outb[0:2]));

	sb_mux_size6_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_1_ccff_tail),
		.mem_out(mem_out[120:122]),
		.mem_outb(mem_outb[120:122]));

	sb_mux_size6_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_2_ccff_tail),
		.mem_out(mem_out[135:137]),
		.mem_outb(mem_outb[135:137]));

	sb_mux_size6_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_3_ccff_tail),
		.mem_out(mem_out[138:140]),
		.mem_outb(mem_outb[138:140]));

	sb_mux_size6_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_4_ccff_tail),
		.mem_out(mem_out[223:225]),
		.mem_outb(mem_outb[223:225]));

	sb_mux_size6_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_15_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_5_ccff_tail),
		.mem_out(mem_out[241:243]),
		.mem_outb(mem_outb[241:243]));

	sb_mux_size6_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_6_ccff_tail),
		.mem_out(mem_out[244:246]),
		.mem_outb(mem_outb[244:246]));

	sb_mux_size6_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_7_ccff_tail),
		.mem_out(mem_out[256:258]),
		.mem_outb(mem_outb[256:258]));

	sb_mux_size5_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_0_ccff_tail),
		.mem_out(mem_out[3:5]),
		.mem_outb(mem_outb[3:5]));

	sb_mux_size5_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_1_ccff_tail),
		.mem_out(mem_out[18:20]),
		.mem_outb(mem_outb[18:20]));

	sb_mux_size5_mem mem_top_track_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_2_ccff_tail),
		.mem_out(mem_out[21:23]),
		.mem_outb(mem_outb[21:23]));

	sb_mux_size5_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_3_ccff_tail),
		.mem_out(mem_out[117:119]),
		.mem_outb(mem_outb[117:119]));

	sb_mux_size5_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_4_ccff_tail),
		.mem_out(mem_out[123:125]),
		.mem_outb(mem_outb[123:125]));

	sb_mux_size5_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_5_ccff_tail),
		.mem_out(mem_out[126:128]),
		.mem_outb(mem_outb[126:128]));

	sb_mux_size5_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_6_ccff_tail),
		.mem_out(mem_out[129:131]),
		.mem_outb(mem_outb[129:131]));

	sb_mux_size5_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_7_ccff_tail),
		.mem_out(mem_out[141:143]),
		.mem_outb(mem_outb[141:143]));

	sb_mux_size5_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_8_ccff_tail),
		.mem_out(mem_out[144:146]),
		.mem_outb(mem_outb[144:146]));

	sb_mux_size5_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_9_ccff_tail),
		.mem_out(mem_out[147:149]),
		.mem_outb(mem_outb[147:149]));

	sb_mux_size5_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_10_ccff_tail),
		.mem_out(mem_out[150:152]),
		.mem_outb(mem_outb[150:152]));

	sb_mux_size5_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_11_ccff_tail),
		.mem_out(mem_out[226:228]),
		.mem_outb(mem_outb[226:228]));

	sb_mux_size5_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_12_ccff_tail),
		.mem_out(mem_out[247:249]),
		.mem_outb(mem_outb[247:249]));

	sb_mux_size5_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_13_ccff_tail),
		.mem_out(mem_out[250:252]),
		.mem_outb(mem_outb[250:252]));

	sb_mux_size5_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_14_ccff_tail),
		.mem_out(mem_out[253:255]),
		.mem_outb(mem_outb[253:255]));

	sb_mux_size5_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_15_ccff_tail),
		.mem_out(mem_out[259:261]),
		.mem_outb(mem_outb[259:261]));

	sb_mux_size5_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_15_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[262:264]),
		.mem_outb(mem_outb[262:264]));

	sb_mux_size4_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_0_ccff_tail),
		.mem_out(mem_out[6:8]),
		.mem_outb(mem_outb[6:8]));

	sb_mux_size4_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_1_ccff_tail),
		.mem_out(mem_out[9:11]),
		.mem_outb(mem_outb[9:11]));

	sb_mux_size4_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_2_ccff_tail),
		.mem_out(mem_out[12:14]),
		.mem_outb(mem_outb[12:14]));

	sb_mux_size4_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_3_ccff_tail),
		.mem_out(mem_out[15:17]),
		.mem_outb(mem_outb[15:17]));

	sb_mux_size4_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_4_ccff_tail),
		.mem_out(mem_out[24:26]),
		.mem_outb(mem_outb[24:26]));

	sb_mux_size4_mem mem_top_track_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_5_ccff_tail),
		.mem_out(mem_out[27:29]),
		.mem_outb(mem_outb[27:29]));

	sb_mux_size4_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_6_ccff_tail),
		.mem_out(mem_out[30:32]),
		.mem_outb(mem_outb[30:32]));

	sb_mux_size4_mem mem_top_track_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_7_ccff_tail),
		.mem_out(mem_out[33:35]),
		.mem_outb(mem_outb[33:35]));

	sb_mux_size4_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_8_ccff_tail),
		.mem_out(mem_out[36:38]),
		.mem_outb(mem_outb[36:38]));

	sb_mux_size4_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_9_ccff_tail),
		.mem_out(mem_out[132:134]),
		.mem_outb(mem_outb[132:134]));

	sb_mux_size4_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_10_ccff_tail),
		.mem_out(mem_out[153:155]),
		.mem_outb(mem_outb[153:155]));

	sb_mux_size4_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_11_ccff_tail),
		.mem_out(mem_out[156:158]),
		.mem_outb(mem_outb[156:158]));

	sb_mux_size4_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_12_ccff_tail),
		.mem_out(mem_out[229:231]),
		.mem_outb(mem_outb[229:231]));

	sb_mux_size4_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_13_ccff_tail),
		.mem_out(mem_out[232:234]),
		.mem_outb(mem_outb[232:234]));

	sb_mux_size4_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_14_ccff_tail),
		.mem_out(mem_out[235:237]),
		.mem_outb(mem_outb[235:237]));

	sb_mux_size4_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_15_ccff_tail),
		.mem_out(mem_out[238:240]),
		.mem_outb(mem_outb[238:240]));

	sb_mux_size3_mem mem_top_track_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[39:40]),
		.mem_outb(mem_outb[39:40]));

	sb_mux_size3_mem mem_top_track_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[41:42]),
		.mem_outb(mem_outb[41:42]));

	sb_mux_size3_mem mem_top_track_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[43:44]),
		.mem_outb(mem_outb[43:44]));

	sb_mux_size3_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[45:46]),
		.mem_outb(mem_outb[45:46]));

	sb_mux_size3_mem mem_top_track_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[47:48]),
		.mem_outb(mem_outb[47:48]));

	sb_mux_size2_mem mem_top_track_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_0_ccff_tail),
		.mem_out(mem_out[49:50]),
		.mem_outb(mem_outb[49:50]));

	sb_mux_size2_mem mem_top_track_62 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_1_ccff_tail),
		.mem_out(mem_out[51:52]),
		.mem_outb(mem_outb[51:52]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[53:54]),
		.mem_outb(mem_outb[53:54]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[55:56]),
		.mem_outb(mem_outb[55:56]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[57:58]),
		.mem_outb(mem_outb[57:58]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[59:60]),
		.mem_outb(mem_outb[59:60]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[61:62]),
		.mem_outb(mem_outb[61:62]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[63:64]),
		.mem_outb(mem_outb[63:64]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[65:66]),
		.mem_outb(mem_outb[65:66]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[67:68]),
		.mem_outb(mem_outb[67:68]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[69:70]),
		.mem_outb(mem_outb[69:70]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[71:72]),
		.mem_outb(mem_outb[71:72]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[73:74]),
		.mem_outb(mem_outb[73:74]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[75:76]),
		.mem_outb(mem_outb[75:76]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[77:78]),
		.mem_outb(mem_outb[77:78]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[79:80]),
		.mem_outb(mem_outb[79:80]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[81:82]),
		.mem_outb(mem_outb[81:82]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[83:84]),
		.mem_outb(mem_outb[83:84]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[85:86]),
		.mem_outb(mem_outb[85:86]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[87:88]),
		.mem_outb(mem_outb[87:88]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[89:90]),
		.mem_outb(mem_outb[89:90]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[91:92]),
		.mem_outb(mem_outb[91:92]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[93:94]),
		.mem_outb(mem_outb[93:94]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[95:96]),
		.mem_outb(mem_outb[95:96]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[97:98]),
		.mem_outb(mem_outb[97:98]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[99:100]),
		.mem_outb(mem_outb[99:100]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[101:102]),
		.mem_outb(mem_outb[101:102]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[103:104]),
		.mem_outb(mem_outb[103:104]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[105:106]),
		.mem_outb(mem_outb[105:106]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[107:108]),
		.mem_outb(mem_outb[107:108]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[109:110]),
		.mem_outb(mem_outb[109:110]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[111:112]),
		.mem_outb(mem_outb[111:112]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[113:114]),
		.mem_outb(mem_outb[113:114]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[115:116]),
		.mem_outb(mem_outb[115:116]));

	clk_mux_size3_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[159:160]),
		.mem_outb(mem_outb[159:160]));

	clk_mux_size3_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[161:162]),
		.mem_outb(mem_outb[161:162]));

	clk_mux_size3_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[163:164]),
		.mem_outb(mem_outb[163:164]));

	clk_mux_size3_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[165:166]),
		.mem_outb(mem_outb[165:166]));

	clk_mux_size3_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[167:168]),
		.mem_outb(mem_outb[167:168]));

	clk_mux_size3_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[169:170]),
		.mem_outb(mem_outb[169:170]));

	clk_mux_size3_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[171:172]),
		.mem_outb(mem_outb[171:172]));

	clk_mux_size3_mem mem_bottom_track_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[173:174]),
		.mem_outb(mem_outb[173:174]));

	clk_mux_size3_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[175:176]),
		.mem_outb(mem_outb[175:176]));

	clk_mux_size3_mem mem_bottom_track_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[177:178]),
		.mem_outb(mem_outb[177:178]));

	clk_mux_size3_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[179:180]),
		.mem_outb(mem_outb[179:180]));

	clk_mux_size3_mem mem_bottom_track_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[181:182]),
		.mem_outb(mem_outb[181:182]));

	clk_mux_size3_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[183:184]),
		.mem_outb(mem_outb[183:184]));

	clk_mux_size3_mem mem_bottom_track_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[185:186]),
		.mem_outb(mem_outb[185:186]));

	clk_mux_size3_mem mem_bottom_track_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[187:188]),
		.mem_outb(mem_outb[187:188]));

	clk_mux_size3_mem mem_bottom_track_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[189:190]),
		.mem_outb(mem_outb[189:190]));

	clk_mux_size3_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[191:192]),
		.mem_outb(mem_outb[191:192]));

	clk_mux_size3_mem mem_bottom_track_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[193:194]),
		.mem_outb(mem_outb[193:194]));

	clk_mux_size3_mem mem_bottom_track_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[195:196]),
		.mem_outb(mem_outb[195:196]));

	clk_mux_size3_mem mem_bottom_track_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[197:198]),
		.mem_outb(mem_outb[197:198]));

	clk_mux_size3_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[199:200]),
		.mem_outb(mem_outb[199:200]));

	clk_mux_size3_mem mem_bottom_track_43 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[201:202]),
		.mem_outb(mem_outb[201:202]));

	clk_mux_size3_mem mem_bottom_track_45 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[203:204]),
		.mem_outb(mem_outb[203:204]));

	clk_mux_size3_mem mem_bottom_track_47 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[205:206]),
		.mem_outb(mem_outb[205:206]));

	clk_mux_size3_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[207:208]),
		.mem_outb(mem_outb[207:208]));

	clk_mux_size3_mem mem_bottom_track_51 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[209:210]),
		.mem_outb(mem_outb[209:210]));

	clk_mux_size3_mem mem_bottom_track_53 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[211:212]),
		.mem_outb(mem_outb[211:212]));

	clk_mux_size3_mem mem_bottom_track_55 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[213:214]),
		.mem_outb(mem_outb[213:214]));

	clk_mux_size3_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[215:216]),
		.mem_outb(mem_outb[215:216]));

	clk_mux_size3_mem mem_bottom_track_59 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[217:218]),
		.mem_outb(mem_outb[217:218]));

	clk_mux_size3_mem mem_bottom_track_61 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[219:220]),
		.mem_outb(mem_outb[219:220]));

	clk_mux_size3_mem mem_bottom_track_63 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[221:222]),
		.mem_outb(mem_outb[221:222]));

endmodule
// ----- END Verilog module for sb_0__config_group_mem_size265 -----




// ----- Verilog module for sb_1__config_group_mem_size344 -----
module sb_1__config_group_mem_size344(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:343] mem_out;
//----- OUTPUT PORTS -----
output [0:343] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size11_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size11_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size11_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[22:25]),
		.mem_outb(mem_outb[22:25]));

	sb_mux_size11_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[26:29]),
		.mem_outb(mem_outb[26:29]));

	sb_mux_size11_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_4_ccff_tail),
		.mem_out(mem_out[140:143]),
		.mem_outb(mem_outb[140:143]));

	sb_mux_size11_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_5_ccff_tail),
		.mem_out(mem_out[144:147]),
		.mem_outb(mem_outb[144:147]));

	sb_mux_size11_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_6_ccff_tail),
		.mem_out(mem_out[148:151]),
		.mem_outb(mem_outb[148:151]));

	sb_mux_size11_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_7_ccff_tail),
		.mem_out(mem_out[172:175]),
		.mem_outb(mem_outb[172:175]));

	sb_mux_size11_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_8_ccff_tail),
		.mem_out(mem_out[176:179]),
		.mem_outb(mem_outb[176:179]));

	sb_mux_size11_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_9_ccff_tail),
		.mem_out(mem_out[194:197]),
		.mem_outb(mem_outb[194:197]));

	sb_mux_size11_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_10_ccff_tail),
		.mem_out(mem_out[198:201]),
		.mem_outb(mem_outb[198:201]));

	sb_mux_size11_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_11_ccff_tail),
		.mem_out(mem_out[312:315]),
		.mem_outb(mem_outb[312:315]));

	sb_mux_size11_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_12_ccff_tail),
		.mem_out(mem_out[316:319]),
		.mem_outb(mem_outb[316:319]));

	sb_mux_size11_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_13_ccff_tail),
		.mem_out(mem_out[320:323]),
		.mem_outb(mem_outb[320:323]));

	sb_mux_size9_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size9_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size9_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_2_ccff_tail),
		.mem_out(mem_out[30:33]),
		.mem_outb(mem_outb[30:33]));

	sb_mux_size9_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_3_ccff_tail),
		.mem_out(mem_out[34:37]),
		.mem_outb(mem_outb[34:37]));

	sb_mux_size9_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_4_ccff_tail),
		.mem_out(mem_out[38:41]),
		.mem_outb(mem_outb[38:41]));

	sb_mux_size9_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_5_ccff_tail),
		.mem_out(mem_out[42:45]),
		.mem_outb(mem_outb[42:45]));

	sb_mux_size9_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_6_ccff_tail),
		.mem_out(mem_out[152:155]),
		.mem_outb(mem_outb[152:155]));

	sb_mux_size9_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_7_ccff_tail),
		.mem_out(mem_out[156:159]),
		.mem_outb(mem_outb[156:159]));

	sb_mux_size9_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_8_ccff_tail),
		.mem_out(mem_out[160:163]),
		.mem_outb(mem_outb[160:163]));

	sb_mux_size9_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_9_ccff_tail),
		.mem_out(mem_out[180:183]),
		.mem_outb(mem_outb[180:183]));

	sb_mux_size9_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_10_ccff_tail),
		.mem_out(mem_out[184:187]),
		.mem_outb(mem_outb[184:187]));

	sb_mux_size9_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_11_ccff_tail),
		.mem_out(mem_out[202:205]),
		.mem_outb(mem_outb[202:205]));

	sb_mux_size9_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_12_ccff_tail),
		.mem_out(mem_out[206:209]),
		.mem_outb(mem_outb[206:209]));

	sb_mux_size9_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_13_ccff_tail),
		.mem_out(mem_out[210:213]),
		.mem_outb(mem_outb[210:213]));

	sb_mux_size9_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_14_ccff_tail),
		.mem_out(mem_out[214:217]),
		.mem_outb(mem_outb[214:217]));

	sb_mux_size9_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_15_ccff_tail),
		.mem_out(mem_out[324:327]),
		.mem_outb(mem_outb[324:327]));

	sb_mux_size9_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_15_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_16_ccff_tail),
		.mem_out(mem_out[328:331]),
		.mem_outb(mem_outb[328:331]));

	sb_mux_size9_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_16_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_17_ccff_tail),
		.mem_out(mem_out[332:335]),
		.mem_outb(mem_outb[332:335]));

	sb_mux_size7_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_0_ccff_tail),
		.mem_out(mem_out[16:18]),
		.mem_outb(mem_outb[16:18]));

	sb_mux_size7_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_1_ccff_tail),
		.mem_out(mem_out[19:21]),
		.mem_outb(mem_outb[19:21]));

	sb_mux_size7_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_2_ccff_tail),
		.mem_out(mem_out[46:48]),
		.mem_outb(mem_outb[46:48]));

	sb_mux_size7_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_3_ccff_tail),
		.mem_out(mem_out[49:51]),
		.mem_outb(mem_outb[49:51]));

	sb_mux_size7_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_4_ccff_tail),
		.mem_out(mem_out[188:190]),
		.mem_outb(mem_outb[188:190]));

	sb_mux_size7_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_5_ccff_tail),
		.mem_out(mem_out[191:193]),
		.mem_outb(mem_outb[191:193]));

	sb_mux_size7_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_6_ccff_tail),
		.mem_out(mem_out[218:220]),
		.mem_outb(mem_outb[218:220]));

	sb_mux_size7_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_7_ccff_tail),
		.mem_out(mem_out[221:223]),
		.mem_outb(mem_outb[221:223]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[52:53]),
		.mem_outb(mem_outb[52:53]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[54:55]),
		.mem_outb(mem_outb[54:55]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[64:65]),
		.mem_outb(mem_outb[64:65]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[66:67]),
		.mem_outb(mem_outb[66:67]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[68:69]),
		.mem_outb(mem_outb[68:69]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[70:71]),
		.mem_outb(mem_outb[70:71]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[72:73]),
		.mem_outb(mem_outb[72:73]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[74:75]),
		.mem_outb(mem_outb[74:75]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[76:77]),
		.mem_outb(mem_outb[76:77]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[78:79]),
		.mem_outb(mem_outb[78:79]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[80:81]),
		.mem_outb(mem_outb[80:81]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[82:83]),
		.mem_outb(mem_outb[82:83]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[84:85]),
		.mem_outb(mem_outb[84:85]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[86:87]),
		.mem_outb(mem_outb[86:87]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[88:89]),
		.mem_outb(mem_outb[88:89]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[94:95]),
		.mem_outb(mem_outb[94:95]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[96:97]),
		.mem_outb(mem_outb[96:97]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[98:99]),
		.mem_outb(mem_outb[98:99]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[224:225]),
		.mem_outb(mem_outb[224:225]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[226:227]),
		.mem_outb(mem_outb[226:227]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[228:229]),
		.mem_outb(mem_outb[228:229]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[230:231]),
		.mem_outb(mem_outb[230:231]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[232:233]),
		.mem_outb(mem_outb[232:233]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[234:235]),
		.mem_outb(mem_outb[234:235]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[236:237]),
		.mem_outb(mem_outb[236:237]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[238:239]),
		.mem_outb(mem_outb[238:239]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[240:241]),
		.mem_outb(mem_outb[240:241]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[242:243]),
		.mem_outb(mem_outb[242:243]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[244:245]),
		.mem_outb(mem_outb[244:245]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[246:247]),
		.mem_outb(mem_outb[246:247]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[248:249]),
		.mem_outb(mem_outb[248:249]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[250:251]),
		.mem_outb(mem_outb[250:251]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[252:253]),
		.mem_outb(mem_outb[252:253]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[254:255]),
		.mem_outb(mem_outb[254:255]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[256:257]),
		.mem_outb(mem_outb[256:257]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[258:259]),
		.mem_outb(mem_outb[258:259]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[260:261]),
		.mem_outb(mem_outb[260:261]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[262:263]),
		.mem_outb(mem_outb[262:263]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[264:265]),
		.mem_outb(mem_outb[264:265]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[266:267]),
		.mem_outb(mem_outb[266:267]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[268:269]),
		.mem_outb(mem_outb[268:269]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[270:271]),
		.mem_outb(mem_outb[270:271]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[272:273]),
		.mem_outb(mem_outb[272:273]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[274:275]),
		.mem_outb(mem_outb[274:275]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[276:277]),
		.mem_outb(mem_outb[276:277]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[278:279]),
		.mem_outb(mem_outb[278:279]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[280:281]),
		.mem_outb(mem_outb[280:281]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[282:283]),
		.mem_outb(mem_outb[282:283]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[284:285]),
		.mem_outb(mem_outb[284:285]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[286:287]),
		.mem_outb(mem_outb[286:287]));

	sb_mux_size10_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[116:119]),
		.mem_outb(mem_outb[116:119]));

	sb_mux_size10_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[120:123]),
		.mem_outb(mem_outb[120:123]));

	sb_mux_size10_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_2_ccff_tail),
		.mem_out(mem_out[124:127]),
		.mem_outb(mem_outb[124:127]));

	sb_mux_size10_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_3_ccff_tail),
		.mem_out(mem_out[128:131]),
		.mem_outb(mem_outb[128:131]));

	sb_mux_size10_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_4_ccff_tail),
		.mem_out(mem_out[288:291]),
		.mem_outb(mem_outb[288:291]));

	sb_mux_size10_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_5_ccff_tail),
		.mem_out(mem_out[292:295]),
		.mem_outb(mem_outb[292:295]));

	sb_mux_size10_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_6_ccff_tail),
		.mem_out(mem_out[296:299]),
		.mem_outb(mem_outb[296:299]));

	sb_mux_size10_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_7_ccff_tail),
		.mem_out(mem_out[300:303]),
		.mem_outb(mem_outb[300:303]));

	sb_mux_size8_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[132:135]),
		.mem_outb(mem_outb[132:135]));

	sb_mux_size8_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[136:139]),
		.mem_outb(mem_outb[136:139]));

	sb_mux_size8_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[164:167]),
		.mem_outb(mem_outb[164:167]));

	sb_mux_size8_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[168:171]),
		.mem_outb(mem_outb[168:171]));

	sb_mux_size8_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[304:307]),
		.mem_outb(mem_outb[304:307]));

	sb_mux_size8_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[308:311]),
		.mem_outb(mem_outb[308:311]));

	sb_mux_size8_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_17_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[336:339]),
		.mem_outb(mem_outb[336:339]));

	sb_mux_size8_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[340:343]),
		.mem_outb(mem_outb[340:343]));

endmodule
// ----- END Verilog module for sb_1__config_group_mem_size344 -----




// ----- Verilog module for sb_2__config_group_mem_size408 -----
module sb_2__config_group_mem_size408(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:407] mem_out;
//----- OUTPUT PORTS -----
output [0:407] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size11_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size11_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size11_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[22:25]),
		.mem_outb(mem_outb[22:25]));

	sb_mux_size11_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[26:29]),
		.mem_outb(mem_outb[26:29]));

	sb_mux_size11_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_4_ccff_tail),
		.mem_out(mem_out[140:143]),
		.mem_outb(mem_outb[140:143]));

	sb_mux_size11_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_5_ccff_tail),
		.mem_out(mem_out[144:147]),
		.mem_outb(mem_outb[144:147]));

	sb_mux_size11_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_6_ccff_tail),
		.mem_out(mem_out[148:151]),
		.mem_outb(mem_outb[148:151]));

	sb_mux_size11_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_7_ccff_tail),
		.mem_out(mem_out[236:239]),
		.mem_outb(mem_outb[236:239]));

	sb_mux_size11_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_8_ccff_tail),
		.mem_out(mem_out[240:243]),
		.mem_outb(mem_outb[240:243]));

	sb_mux_size11_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_9_ccff_tail),
		.mem_out(mem_out[258:261]),
		.mem_outb(mem_outb[258:261]));

	sb_mux_size11_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_10_ccff_tail),
		.mem_out(mem_out[262:265]),
		.mem_outb(mem_outb[262:265]));

	sb_mux_size11_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_11_ccff_tail),
		.mem_out(mem_out[376:379]),
		.mem_outb(mem_outb[376:379]));

	sb_mux_size11_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_12_ccff_tail),
		.mem_out(mem_out[380:383]),
		.mem_outb(mem_outb[380:383]));

	sb_mux_size11_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_13_ccff_tail),
		.mem_out(mem_out[384:387]),
		.mem_outb(mem_outb[384:387]));

	sb_mux_size9_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size9_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size9_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_2_ccff_tail),
		.mem_out(mem_out[30:33]),
		.mem_outb(mem_outb[30:33]));

	sb_mux_size9_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_3_ccff_tail),
		.mem_out(mem_out[34:37]),
		.mem_outb(mem_outb[34:37]));

	sb_mux_size9_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_4_ccff_tail),
		.mem_out(mem_out[38:41]),
		.mem_outb(mem_outb[38:41]));

	sb_mux_size9_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_5_ccff_tail),
		.mem_out(mem_out[42:45]),
		.mem_outb(mem_outb[42:45]));

	sb_mux_size9_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_6_ccff_tail),
		.mem_out(mem_out[152:155]),
		.mem_outb(mem_outb[152:155]));

	sb_mux_size9_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_7_ccff_tail),
		.mem_out(mem_out[156:159]),
		.mem_outb(mem_outb[156:159]));

	sb_mux_size9_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_8_ccff_tail),
		.mem_out(mem_out[160:163]),
		.mem_outb(mem_outb[160:163]));

	sb_mux_size9_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_9_ccff_tail),
		.mem_out(mem_out[244:247]),
		.mem_outb(mem_outb[244:247]));

	sb_mux_size9_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_10_ccff_tail),
		.mem_out(mem_out[248:251]),
		.mem_outb(mem_outb[248:251]));

	sb_mux_size9_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_11_ccff_tail),
		.mem_out(mem_out[266:269]),
		.mem_outb(mem_outb[266:269]));

	sb_mux_size9_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_12_ccff_tail),
		.mem_out(mem_out[270:273]),
		.mem_outb(mem_outb[270:273]));

	sb_mux_size9_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_13_ccff_tail),
		.mem_out(mem_out[274:277]),
		.mem_outb(mem_outb[274:277]));

	sb_mux_size9_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_14_ccff_tail),
		.mem_out(mem_out[278:281]),
		.mem_outb(mem_outb[278:281]));

	sb_mux_size9_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_15_ccff_tail),
		.mem_out(mem_out[388:391]),
		.mem_outb(mem_outb[388:391]));

	sb_mux_size9_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_15_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_16_ccff_tail),
		.mem_out(mem_out[392:395]),
		.mem_outb(mem_outb[392:395]));

	sb_mux_size9_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_16_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_17_ccff_tail),
		.mem_out(mem_out[396:399]),
		.mem_outb(mem_outb[396:399]));

	sb_mux_size7_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_0_ccff_tail),
		.mem_out(mem_out[16:18]),
		.mem_outb(mem_outb[16:18]));

	sb_mux_size7_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_1_ccff_tail),
		.mem_out(mem_out[19:21]),
		.mem_outb(mem_outb[19:21]));

	sb_mux_size7_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_2_ccff_tail),
		.mem_out(mem_out[46:48]),
		.mem_outb(mem_outb[46:48]));

	sb_mux_size7_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_3_ccff_tail),
		.mem_out(mem_out[49:51]),
		.mem_outb(mem_outb[49:51]));

	sb_mux_size7_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_4_ccff_tail),
		.mem_out(mem_out[252:254]),
		.mem_outb(mem_outb[252:254]));

	sb_mux_size7_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_5_ccff_tail),
		.mem_out(mem_out[255:257]),
		.mem_outb(mem_outb[255:257]));

	sb_mux_size7_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_6_ccff_tail),
		.mem_out(mem_out[282:284]),
		.mem_outb(mem_outb[282:284]));

	sb_mux_size7_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_7_ccff_tail),
		.mem_out(mem_out[285:287]),
		.mem_outb(mem_outb[285:287]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[52:53]),
		.mem_outb(mem_outb[52:53]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[54:55]),
		.mem_outb(mem_outb[54:55]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[64:65]),
		.mem_outb(mem_outb[64:65]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[66:67]),
		.mem_outb(mem_outb[66:67]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[68:69]),
		.mem_outb(mem_outb[68:69]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[70:71]),
		.mem_outb(mem_outb[70:71]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[72:73]),
		.mem_outb(mem_outb[72:73]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[74:75]),
		.mem_outb(mem_outb[74:75]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[76:77]),
		.mem_outb(mem_outb[76:77]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[78:79]),
		.mem_outb(mem_outb[78:79]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[80:81]),
		.mem_outb(mem_outb[80:81]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[82:83]),
		.mem_outb(mem_outb[82:83]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[84:85]),
		.mem_outb(mem_outb[84:85]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[86:87]),
		.mem_outb(mem_outb[86:87]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[88:89]),
		.mem_outb(mem_outb[88:89]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[94:95]),
		.mem_outb(mem_outb[94:95]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[96:97]),
		.mem_outb(mem_outb[96:97]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[98:99]),
		.mem_outb(mem_outb[98:99]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	clk_mux_size3_mem mem_right_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[172:173]),
		.mem_outb(mem_outb[172:173]));

	clk_mux_size3_mem mem_right_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[174:175]),
		.mem_outb(mem_outb[174:175]));

	clk_mux_size3_mem mem_right_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[176:177]),
		.mem_outb(mem_outb[176:177]));

	clk_mux_size3_mem mem_right_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[178:179]),
		.mem_outb(mem_outb[178:179]));

	clk_mux_size3_mem mem_right_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[180:181]),
		.mem_outb(mem_outb[180:181]));

	clk_mux_size3_mem mem_right_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[182:183]),
		.mem_outb(mem_outb[182:183]));

	clk_mux_size3_mem mem_right_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[184:185]),
		.mem_outb(mem_outb[184:185]));

	clk_mux_size3_mem mem_right_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[186:187]),
		.mem_outb(mem_outb[186:187]));

	clk_mux_size3_mem mem_right_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[188:189]),
		.mem_outb(mem_outb[188:189]));

	clk_mux_size3_mem mem_right_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[190:191]),
		.mem_outb(mem_outb[190:191]));

	clk_mux_size3_mem mem_right_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[192:193]),
		.mem_outb(mem_outb[192:193]));

	clk_mux_size3_mem mem_right_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[194:195]),
		.mem_outb(mem_outb[194:195]));

	clk_mux_size3_mem mem_right_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[196:197]),
		.mem_outb(mem_outb[196:197]));

	clk_mux_size3_mem mem_right_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[198:199]),
		.mem_outb(mem_outb[198:199]));

	clk_mux_size3_mem mem_right_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[200:201]),
		.mem_outb(mem_outb[200:201]));

	clk_mux_size3_mem mem_right_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[202:203]),
		.mem_outb(mem_outb[202:203]));

	clk_mux_size3_mem mem_right_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[204:205]),
		.mem_outb(mem_outb[204:205]));

	clk_mux_size3_mem mem_right_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[206:207]),
		.mem_outb(mem_outb[206:207]));

	clk_mux_size3_mem mem_right_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[208:209]),
		.mem_outb(mem_outb[208:209]));

	clk_mux_size3_mem mem_right_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[210:211]),
		.mem_outb(mem_outb[210:211]));

	clk_mux_size3_mem mem_right_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[212:213]),
		.mem_outb(mem_outb[212:213]));

	clk_mux_size3_mem mem_right_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[214:215]),
		.mem_outb(mem_outb[214:215]));

	clk_mux_size3_mem mem_right_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[216:217]),
		.mem_outb(mem_outb[216:217]));

	clk_mux_size3_mem mem_right_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[218:219]),
		.mem_outb(mem_outb[218:219]));

	clk_mux_size3_mem mem_right_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[220:221]),
		.mem_outb(mem_outb[220:221]));

	clk_mux_size3_mem mem_right_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[222:223]),
		.mem_outb(mem_outb[222:223]));

	clk_mux_size3_mem mem_right_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[224:225]),
		.mem_outb(mem_outb[224:225]));

	clk_mux_size3_mem mem_right_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[226:227]),
		.mem_outb(mem_outb[226:227]));

	clk_mux_size3_mem mem_right_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[228:229]),
		.mem_outb(mem_outb[228:229]));

	clk_mux_size3_mem mem_right_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[230:231]),
		.mem_outb(mem_outb[230:231]));

	clk_mux_size3_mem mem_right_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[232:233]),
		.mem_outb(mem_outb[232:233]));

	clk_mux_size3_mem mem_right_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[234:235]),
		.mem_outb(mem_outb[234:235]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_64_ccff_tail),
		.mem_out(mem_out[288:289]),
		.mem_outb(mem_outb[288:289]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_64_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_65_ccff_tail),
		.mem_out(mem_out[290:291]),
		.mem_outb(mem_outb[290:291]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_65_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_66_ccff_tail),
		.mem_out(mem_out[292:293]),
		.mem_outb(mem_outb[292:293]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_66_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_67_ccff_tail),
		.mem_out(mem_out[294:295]),
		.mem_outb(mem_outb[294:295]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_67_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_68_ccff_tail),
		.mem_out(mem_out[296:297]),
		.mem_outb(mem_outb[296:297]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_68_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_69_ccff_tail),
		.mem_out(mem_out[298:299]),
		.mem_outb(mem_outb[298:299]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_69_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_70_ccff_tail),
		.mem_out(mem_out[300:301]),
		.mem_outb(mem_outb[300:301]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_70_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_71_ccff_tail),
		.mem_out(mem_out[302:303]),
		.mem_outb(mem_outb[302:303]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_71_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_72_ccff_tail),
		.mem_out(mem_out[304:305]),
		.mem_outb(mem_outb[304:305]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_72_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_73_ccff_tail),
		.mem_out(mem_out[306:307]),
		.mem_outb(mem_outb[306:307]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_73_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_74_ccff_tail),
		.mem_out(mem_out[308:309]),
		.mem_outb(mem_outb[308:309]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_74_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_75_ccff_tail),
		.mem_out(mem_out[310:311]),
		.mem_outb(mem_outb[310:311]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_75_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_76_ccff_tail),
		.mem_out(mem_out[312:313]),
		.mem_outb(mem_outb[312:313]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_76_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_77_ccff_tail),
		.mem_out(mem_out[314:315]),
		.mem_outb(mem_outb[314:315]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_77_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_78_ccff_tail),
		.mem_out(mem_out[316:317]),
		.mem_outb(mem_outb[316:317]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_78_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_79_ccff_tail),
		.mem_out(mem_out[318:319]),
		.mem_outb(mem_outb[318:319]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_79_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_80_ccff_tail),
		.mem_out(mem_out[320:321]),
		.mem_outb(mem_outb[320:321]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_80_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_81_ccff_tail),
		.mem_out(mem_out[322:323]),
		.mem_outb(mem_outb[322:323]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_81_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_82_ccff_tail),
		.mem_out(mem_out[324:325]),
		.mem_outb(mem_outb[324:325]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_82_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_83_ccff_tail),
		.mem_out(mem_out[326:327]),
		.mem_outb(mem_outb[326:327]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_83_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_84_ccff_tail),
		.mem_out(mem_out[328:329]),
		.mem_outb(mem_outb[328:329]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_84_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_85_ccff_tail),
		.mem_out(mem_out[330:331]),
		.mem_outb(mem_outb[330:331]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_85_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_86_ccff_tail),
		.mem_out(mem_out[332:333]),
		.mem_outb(mem_outb[332:333]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_86_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_87_ccff_tail),
		.mem_out(mem_out[334:335]),
		.mem_outb(mem_outb[334:335]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_87_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_88_ccff_tail),
		.mem_out(mem_out[336:337]),
		.mem_outb(mem_outb[336:337]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_88_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_89_ccff_tail),
		.mem_out(mem_out[338:339]),
		.mem_outb(mem_outb[338:339]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_89_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_90_ccff_tail),
		.mem_out(mem_out[340:341]),
		.mem_outb(mem_outb[340:341]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_90_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_91_ccff_tail),
		.mem_out(mem_out[342:343]),
		.mem_outb(mem_outb[342:343]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_91_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_92_ccff_tail),
		.mem_out(mem_out[344:345]),
		.mem_outb(mem_outb[344:345]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_92_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_93_ccff_tail),
		.mem_out(mem_out[346:347]),
		.mem_outb(mem_outb[346:347]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_93_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_94_ccff_tail),
		.mem_out(mem_out[348:349]),
		.mem_outb(mem_outb[348:349]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_94_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_95_ccff_tail),
		.mem_out(mem_out[350:351]),
		.mem_outb(mem_outb[350:351]));

	sb_mux_size10_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[116:119]),
		.mem_outb(mem_outb[116:119]));

	sb_mux_size10_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[120:123]),
		.mem_outb(mem_outb[120:123]));

	sb_mux_size10_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_2_ccff_tail),
		.mem_out(mem_out[124:127]),
		.mem_outb(mem_outb[124:127]));

	sb_mux_size10_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_3_ccff_tail),
		.mem_out(mem_out[128:131]),
		.mem_outb(mem_outb[128:131]));

	sb_mux_size10_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_95_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_4_ccff_tail),
		.mem_out(mem_out[352:355]),
		.mem_outb(mem_outb[352:355]));

	sb_mux_size10_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_5_ccff_tail),
		.mem_out(mem_out[356:359]),
		.mem_outb(mem_outb[356:359]));

	sb_mux_size10_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_6_ccff_tail),
		.mem_out(mem_out[360:363]),
		.mem_outb(mem_outb[360:363]));

	sb_mux_size10_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_7_ccff_tail),
		.mem_out(mem_out[364:367]),
		.mem_outb(mem_outb[364:367]));

	sb_mux_size8_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[132:135]),
		.mem_outb(mem_outb[132:135]));

	sb_mux_size8_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[136:139]),
		.mem_outb(mem_outb[136:139]));

	sb_mux_size8_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[164:167]),
		.mem_outb(mem_outb[164:167]));

	sb_mux_size8_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[168:171]),
		.mem_outb(mem_outb[168:171]));

	sb_mux_size8_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[368:371]),
		.mem_outb(mem_outb[368:371]));

	sb_mux_size8_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[372:375]),
		.mem_outb(mem_outb[372:375]));

	sb_mux_size8_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_17_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[400:403]),
		.mem_outb(mem_outb[400:403]));

	sb_mux_size8_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[404:407]),
		.mem_outb(mem_outb[404:407]));

endmodule
// ----- END Verilog module for sb_2__config_group_mem_size408 -----




// ----- Verilog module for sb_3__config_group_mem_size344 -----
module sb_3__config_group_mem_size344(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:343] mem_out;
//----- OUTPUT PORTS -----
output [0:343] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size11_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size11_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size11_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[22:25]),
		.mem_outb(mem_outb[22:25]));

	sb_mux_size11_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[26:29]),
		.mem_outb(mem_outb[26:29]));

	sb_mux_size11_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_4_ccff_tail),
		.mem_out(mem_out[140:143]),
		.mem_outb(mem_outb[140:143]));

	sb_mux_size11_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_5_ccff_tail),
		.mem_out(mem_out[144:147]),
		.mem_outb(mem_outb[144:147]));

	sb_mux_size11_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_6_ccff_tail),
		.mem_out(mem_out[148:151]),
		.mem_outb(mem_outb[148:151]));

	sb_mux_size11_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_7_ccff_tail),
		.mem_out(mem_out[172:175]),
		.mem_outb(mem_outb[172:175]));

	sb_mux_size11_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_8_ccff_tail),
		.mem_out(mem_out[176:179]),
		.mem_outb(mem_outb[176:179]));

	sb_mux_size11_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_9_ccff_tail),
		.mem_out(mem_out[194:197]),
		.mem_outb(mem_outb[194:197]));

	sb_mux_size11_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_10_ccff_tail),
		.mem_out(mem_out[198:201]),
		.mem_outb(mem_outb[198:201]));

	sb_mux_size11_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_11_ccff_tail),
		.mem_out(mem_out[312:315]),
		.mem_outb(mem_outb[312:315]));

	sb_mux_size11_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_12_ccff_tail),
		.mem_out(mem_out[316:319]),
		.mem_outb(mem_outb[316:319]));

	sb_mux_size11_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_13_ccff_tail),
		.mem_out(mem_out[320:323]),
		.mem_outb(mem_outb[320:323]));

	sb_mux_size9_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size9_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size9_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_2_ccff_tail),
		.mem_out(mem_out[30:33]),
		.mem_outb(mem_outb[30:33]));

	sb_mux_size9_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_3_ccff_tail),
		.mem_out(mem_out[34:37]),
		.mem_outb(mem_outb[34:37]));

	sb_mux_size9_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_4_ccff_tail),
		.mem_out(mem_out[38:41]),
		.mem_outb(mem_outb[38:41]));

	sb_mux_size9_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_5_ccff_tail),
		.mem_out(mem_out[42:45]),
		.mem_outb(mem_outb[42:45]));

	sb_mux_size9_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_6_ccff_tail),
		.mem_out(mem_out[152:155]),
		.mem_outb(mem_outb[152:155]));

	sb_mux_size9_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_7_ccff_tail),
		.mem_out(mem_out[156:159]),
		.mem_outb(mem_outb[156:159]));

	sb_mux_size9_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_8_ccff_tail),
		.mem_out(mem_out[160:163]),
		.mem_outb(mem_outb[160:163]));

	sb_mux_size9_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_9_ccff_tail),
		.mem_out(mem_out[180:183]),
		.mem_outb(mem_outb[180:183]));

	sb_mux_size9_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_10_ccff_tail),
		.mem_out(mem_out[184:187]),
		.mem_outb(mem_outb[184:187]));

	sb_mux_size9_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_11_ccff_tail),
		.mem_out(mem_out[202:205]),
		.mem_outb(mem_outb[202:205]));

	sb_mux_size9_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_12_ccff_tail),
		.mem_out(mem_out[206:209]),
		.mem_outb(mem_outb[206:209]));

	sb_mux_size9_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_13_ccff_tail),
		.mem_out(mem_out[210:213]),
		.mem_outb(mem_outb[210:213]));

	sb_mux_size9_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_14_ccff_tail),
		.mem_out(mem_out[214:217]),
		.mem_outb(mem_outb[214:217]));

	sb_mux_size9_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_15_ccff_tail),
		.mem_out(mem_out[324:327]),
		.mem_outb(mem_outb[324:327]));

	sb_mux_size9_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_15_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_16_ccff_tail),
		.mem_out(mem_out[328:331]),
		.mem_outb(mem_outb[328:331]));

	sb_mux_size9_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_16_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_17_ccff_tail),
		.mem_out(mem_out[332:335]),
		.mem_outb(mem_outb[332:335]));

	sb_mux_size7_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_0_ccff_tail),
		.mem_out(mem_out[16:18]),
		.mem_outb(mem_outb[16:18]));

	sb_mux_size7_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_1_ccff_tail),
		.mem_out(mem_out[19:21]),
		.mem_outb(mem_outb[19:21]));

	sb_mux_size7_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_2_ccff_tail),
		.mem_out(mem_out[46:48]),
		.mem_outb(mem_outb[46:48]));

	sb_mux_size7_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_3_ccff_tail),
		.mem_out(mem_out[49:51]),
		.mem_outb(mem_outb[49:51]));

	sb_mux_size7_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_4_ccff_tail),
		.mem_out(mem_out[188:190]),
		.mem_outb(mem_outb[188:190]));

	sb_mux_size7_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_5_ccff_tail),
		.mem_out(mem_out[191:193]),
		.mem_outb(mem_outb[191:193]));

	sb_mux_size7_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_6_ccff_tail),
		.mem_out(mem_out[218:220]),
		.mem_outb(mem_outb[218:220]));

	sb_mux_size7_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_7_ccff_tail),
		.mem_out(mem_out[221:223]),
		.mem_outb(mem_outb[221:223]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[52:53]),
		.mem_outb(mem_outb[52:53]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[54:55]),
		.mem_outb(mem_outb[54:55]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[64:65]),
		.mem_outb(mem_outb[64:65]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[66:67]),
		.mem_outb(mem_outb[66:67]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[68:69]),
		.mem_outb(mem_outb[68:69]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[70:71]),
		.mem_outb(mem_outb[70:71]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[72:73]),
		.mem_outb(mem_outb[72:73]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[74:75]),
		.mem_outb(mem_outb[74:75]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[76:77]),
		.mem_outb(mem_outb[76:77]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[78:79]),
		.mem_outb(mem_outb[78:79]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[80:81]),
		.mem_outb(mem_outb[80:81]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[82:83]),
		.mem_outb(mem_outb[82:83]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[84:85]),
		.mem_outb(mem_outb[84:85]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[86:87]),
		.mem_outb(mem_outb[86:87]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[88:89]),
		.mem_outb(mem_outb[88:89]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[94:95]),
		.mem_outb(mem_outb[94:95]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[96:97]),
		.mem_outb(mem_outb[96:97]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[98:99]),
		.mem_outb(mem_outb[98:99]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[224:225]),
		.mem_outb(mem_outb[224:225]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[226:227]),
		.mem_outb(mem_outb[226:227]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[228:229]),
		.mem_outb(mem_outb[228:229]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[230:231]),
		.mem_outb(mem_outb[230:231]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[232:233]),
		.mem_outb(mem_outb[232:233]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[234:235]),
		.mem_outb(mem_outb[234:235]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[236:237]),
		.mem_outb(mem_outb[236:237]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[238:239]),
		.mem_outb(mem_outb[238:239]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[240:241]),
		.mem_outb(mem_outb[240:241]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[242:243]),
		.mem_outb(mem_outb[242:243]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[244:245]),
		.mem_outb(mem_outb[244:245]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[246:247]),
		.mem_outb(mem_outb[246:247]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[248:249]),
		.mem_outb(mem_outb[248:249]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[250:251]),
		.mem_outb(mem_outb[250:251]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[252:253]),
		.mem_outb(mem_outb[252:253]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[254:255]),
		.mem_outb(mem_outb[254:255]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[256:257]),
		.mem_outb(mem_outb[256:257]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[258:259]),
		.mem_outb(mem_outb[258:259]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[260:261]),
		.mem_outb(mem_outb[260:261]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[262:263]),
		.mem_outb(mem_outb[262:263]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[264:265]),
		.mem_outb(mem_outb[264:265]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[266:267]),
		.mem_outb(mem_outb[266:267]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[268:269]),
		.mem_outb(mem_outb[268:269]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[270:271]),
		.mem_outb(mem_outb[270:271]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[272:273]),
		.mem_outb(mem_outb[272:273]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[274:275]),
		.mem_outb(mem_outb[274:275]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[276:277]),
		.mem_outb(mem_outb[276:277]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[278:279]),
		.mem_outb(mem_outb[278:279]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[280:281]),
		.mem_outb(mem_outb[280:281]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[282:283]),
		.mem_outb(mem_outb[282:283]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[284:285]),
		.mem_outb(mem_outb[284:285]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[286:287]),
		.mem_outb(mem_outb[286:287]));

	sb_mux_size10_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[116:119]),
		.mem_outb(mem_outb[116:119]));

	sb_mux_size10_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[120:123]),
		.mem_outb(mem_outb[120:123]));

	sb_mux_size10_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_2_ccff_tail),
		.mem_out(mem_out[124:127]),
		.mem_outb(mem_outb[124:127]));

	sb_mux_size10_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_3_ccff_tail),
		.mem_out(mem_out[128:131]),
		.mem_outb(mem_outb[128:131]));

	sb_mux_size10_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_4_ccff_tail),
		.mem_out(mem_out[288:291]),
		.mem_outb(mem_outb[288:291]));

	sb_mux_size10_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_5_ccff_tail),
		.mem_out(mem_out[292:295]),
		.mem_outb(mem_outb[292:295]));

	sb_mux_size10_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_6_ccff_tail),
		.mem_out(mem_out[296:299]),
		.mem_outb(mem_outb[296:299]));

	sb_mux_size10_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_7_ccff_tail),
		.mem_out(mem_out[300:303]),
		.mem_outb(mem_outb[300:303]));

	sb_mux_size8_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[132:135]),
		.mem_outb(mem_outb[132:135]));

	sb_mux_size8_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[136:139]),
		.mem_outb(mem_outb[136:139]));

	sb_mux_size8_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[164:167]),
		.mem_outb(mem_outb[164:167]));

	sb_mux_size8_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[168:171]),
		.mem_outb(mem_outb[168:171]));

	sb_mux_size8_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[304:307]),
		.mem_outb(mem_outb[304:307]));

	sb_mux_size8_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[308:311]),
		.mem_outb(mem_outb[308:311]));

	sb_mux_size8_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_17_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[336:339]),
		.mem_outb(mem_outb[336:339]));

	sb_mux_size8_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[340:343]),
		.mem_outb(mem_outb[340:343]));

endmodule
// ----- END Verilog module for sb_3__config_group_mem_size344 -----




// ----- Verilog module for sb_4__config_group_mem_size244 -----
module sb_4__config_group_mem_size244(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:243] mem_out;
//----- OUTPUT PORTS -----
output [0:243] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	clk_mux_size3_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[0:1]),
		.mem_outb(mem_outb[0:1]));

	clk_mux_size3_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[2:3]),
		.mem_outb(mem_outb[2:3]));

	clk_mux_size3_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[4:5]),
		.mem_outb(mem_outb[4:5]));

	clk_mux_size3_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[6:7]),
		.mem_outb(mem_outb[6:7]));

	clk_mux_size3_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[8:9]),
		.mem_outb(mem_outb[8:9]));

	clk_mux_size3_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[10:11]),
		.mem_outb(mem_outb[10:11]));

	clk_mux_size3_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[12:13]),
		.mem_outb(mem_outb[12:13]));

	clk_mux_size3_mem mem_top_track_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[14:15]),
		.mem_outb(mem_outb[14:15]));

	clk_mux_size3_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[16:17]),
		.mem_outb(mem_outb[16:17]));

	clk_mux_size3_mem mem_top_track_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[18:19]),
		.mem_outb(mem_outb[18:19]));

	clk_mux_size3_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[20:21]),
		.mem_outb(mem_outb[20:21]));

	clk_mux_size3_mem mem_top_track_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[22:23]),
		.mem_outb(mem_outb[22:23]));

	clk_mux_size3_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[24:25]),
		.mem_outb(mem_outb[24:25]));

	clk_mux_size3_mem mem_top_track_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[26:27]),
		.mem_outb(mem_outb[26:27]));

	clk_mux_size3_mem mem_top_track_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[28:29]),
		.mem_outb(mem_outb[28:29]));

	clk_mux_size3_mem mem_top_track_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[30:31]),
		.mem_outb(mem_outb[30:31]));

	clk_mux_size3_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[32:33]),
		.mem_outb(mem_outb[32:33]));

	clk_mux_size3_mem mem_top_track_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[34:35]),
		.mem_outb(mem_outb[34:35]));

	clk_mux_size3_mem mem_top_track_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[36:37]),
		.mem_outb(mem_outb[36:37]));

	clk_mux_size3_mem mem_top_track_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[38:39]),
		.mem_outb(mem_outb[38:39]));

	clk_mux_size3_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[40:41]),
		.mem_outb(mem_outb[40:41]));

	clk_mux_size3_mem mem_top_track_42 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[42:43]),
		.mem_outb(mem_outb[42:43]));

	clk_mux_size3_mem mem_top_track_44 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[44:45]),
		.mem_outb(mem_outb[44:45]));

	clk_mux_size3_mem mem_top_track_46 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[46:47]),
		.mem_outb(mem_outb[46:47]));

	clk_mux_size3_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[48:49]),
		.mem_outb(mem_outb[48:49]));

	clk_mux_size3_mem mem_top_track_50 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[50:51]),
		.mem_outb(mem_outb[50:51]));

	clk_mux_size3_mem mem_top_track_52 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[52:53]),
		.mem_outb(mem_outb[52:53]));

	clk_mux_size3_mem mem_top_track_54 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[54:55]),
		.mem_outb(mem_outb[54:55]));

	clk_mux_size3_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_58 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_60 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_62 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[180:181]),
		.mem_outb(mem_outb[180:181]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[182:183]),
		.mem_outb(mem_outb[182:183]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[184:185]),
		.mem_outb(mem_outb[184:185]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[186:187]),
		.mem_outb(mem_outb[186:187]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[188:189]),
		.mem_outb(mem_outb[188:189]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[190:191]),
		.mem_outb(mem_outb[190:191]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[192:193]),
		.mem_outb(mem_outb[192:193]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[194:195]),
		.mem_outb(mem_outb[194:195]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[196:197]),
		.mem_outb(mem_outb[196:197]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[198:199]),
		.mem_outb(mem_outb[198:199]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[200:201]),
		.mem_outb(mem_outb[200:201]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[202:203]),
		.mem_outb(mem_outb[202:203]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[204:205]),
		.mem_outb(mem_outb[204:205]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[206:207]),
		.mem_outb(mem_outb[206:207]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[208:209]),
		.mem_outb(mem_outb[208:209]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[210:211]),
		.mem_outb(mem_outb[210:211]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[212:213]),
		.mem_outb(mem_outb[212:213]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[214:215]),
		.mem_outb(mem_outb[214:215]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[216:217]),
		.mem_outb(mem_outb[216:217]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[218:219]),
		.mem_outb(mem_outb[218:219]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[220:221]),
		.mem_outb(mem_outb[220:221]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[222:223]),
		.mem_outb(mem_outb[222:223]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[224:225]),
		.mem_outb(mem_outb[224:225]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[226:227]),
		.mem_outb(mem_outb[226:227]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[228:229]),
		.mem_outb(mem_outb[228:229]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[230:231]),
		.mem_outb(mem_outb[230:231]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[232:233]),
		.mem_outb(mem_outb[232:233]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[234:235]),
		.mem_outb(mem_outb[234:235]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[236:237]),
		.mem_outb(mem_outb[236:237]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[238:239]),
		.mem_outb(mem_outb[238:239]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[240:241]),
		.mem_outb(mem_outb[240:241]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[242:243]),
		.mem_outb(mem_outb[242:243]));

	sb_mux_size6_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_0_ccff_tail),
		.mem_out(mem_out[64:66]),
		.mem_outb(mem_outb[64:66]));

	sb_mux_size6_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_1_ccff_tail),
		.mem_out(mem_out[67:69]),
		.mem_outb(mem_outb[67:69]));

	sb_mux_size6_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_2_ccff_tail),
		.mem_out(mem_out[82:84]),
		.mem_outb(mem_outb[82:84]));

	sb_mux_size6_mem mem_right_track_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_3_ccff_tail),
		.mem_out(mem_out[85:87]),
		.mem_outb(mem_outb[85:87]));

	sb_mux_size5_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_0_ccff_tail),
		.mem_out(mem_out[70:72]),
		.mem_outb(mem_outb[70:72]));

	sb_mux_size5_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_1_ccff_tail),
		.mem_out(mem_out[73:75]),
		.mem_outb(mem_outb[73:75]));

	sb_mux_size5_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_2_ccff_tail),
		.mem_out(mem_out[76:78]),
		.mem_outb(mem_outb[76:78]));

	sb_mux_size5_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_3_ccff_tail),
		.mem_out(mem_out[79:81]),
		.mem_outb(mem_outb[79:81]));

	sb_mux_size5_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_4_ccff_tail),
		.mem_out(mem_out[88:90]),
		.mem_outb(mem_outb[88:90]));

	sb_mux_size5_mem mem_right_track_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_5_ccff_tail),
		.mem_out(mem_out[91:93]),
		.mem_outb(mem_outb[91:93]));

	sb_mux_size5_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_6_ccff_tail),
		.mem_out(mem_out[94:96]),
		.mem_outb(mem_outb[94:96]));

	sb_mux_size5_mem mem_right_track_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_7_ccff_tail),
		.mem_out(mem_out[97:99]),
		.mem_outb(mem_outb[97:99]));

	sb_mux_size3_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	sb_mux_size3_mem mem_right_track_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	sb_mux_size3_mem mem_right_track_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	sb_mux_size3_mem mem_right_track_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	sb_mux_size3_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	sb_mux_size3_mem mem_right_track_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	sb_mux_size3_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[140:141]),
		.mem_outb(mem_outb[140:141]));

	sb_mux_size3_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[142:143]),
		.mem_outb(mem_outb[142:143]));

	sb_mux_size3_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_17_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[152:153]),
		.mem_outb(mem_outb[152:153]));

	sb_mux_size3_mem mem_bottom_track_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[154:155]),
		.mem_outb(mem_outb[154:155]));

	sb_mux_size2_mem mem_right_track_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_0_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	sb_mux_size2_mem mem_right_track_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_1_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	sb_mux_size2_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_2_ccff_tail),
		.mem_out(mem_out[116:117]),
		.mem_outb(mem_outb[116:117]));

	sb_mux_size2_mem mem_right_track_42 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_3_ccff_tail),
		.mem_out(mem_out[118:119]),
		.mem_outb(mem_outb[118:119]));

	sb_mux_size2_mem mem_right_track_44 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_4_ccff_tail),
		.mem_out(mem_out[120:121]),
		.mem_outb(mem_outb[120:121]));

	sb_mux_size2_mem mem_right_track_46 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_5_ccff_tail),
		.mem_out(mem_out[122:123]),
		.mem_outb(mem_outb[122:123]));

	sb_mux_size2_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_6_ccff_tail),
		.mem_out(mem_out[124:125]),
		.mem_outb(mem_outb[124:125]));

	sb_mux_size2_mem mem_right_track_50 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_7_ccff_tail),
		.mem_out(mem_out[126:127]),
		.mem_outb(mem_outb[126:127]));

	sb_mux_size2_mem mem_right_track_52 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_8_ccff_tail),
		.mem_out(mem_out[128:129]),
		.mem_outb(mem_outb[128:129]));

	sb_mux_size2_mem mem_right_track_54 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_9_ccff_tail),
		.mem_out(mem_out[130:131]),
		.mem_outb(mem_outb[130:131]));

	sb_mux_size2_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_10_ccff_tail),
		.mem_out(mem_out[132:133]),
		.mem_outb(mem_outb[132:133]));

	sb_mux_size2_mem mem_right_track_58 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_11_ccff_tail),
		.mem_out(mem_out[134:135]),
		.mem_outb(mem_outb[134:135]));

	sb_mux_size2_mem mem_right_track_60 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_12_ccff_tail),
		.mem_out(mem_out[136:137]),
		.mem_outb(mem_outb[136:137]));

	sb_mux_size2_mem mem_right_track_62 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_13_ccff_tail),
		.mem_out(mem_out[138:139]),
		.mem_outb(mem_outb[138:139]));

	sb_mux_size2_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_14_ccff_tail),
		.mem_out(mem_out[144:145]),
		.mem_outb(mem_outb[144:145]));

	sb_mux_size2_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_15_ccff_tail),
		.mem_out(mem_out[146:147]),
		.mem_outb(mem_outb[146:147]));

	sb_mux_size2_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_15_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_16_ccff_tail),
		.mem_out(mem_out[148:149]),
		.mem_outb(mem_outb[148:149]));

	sb_mux_size2_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_16_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_17_ccff_tail),
		.mem_out(mem_out[150:151]),
		.mem_outb(mem_outb[150:151]));

	sb_mux_size2_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size3_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_18_ccff_tail),
		.mem_out(mem_out[156:157]),
		.mem_outb(mem_outb[156:157]));

	sb_mux_size2_mem mem_bottom_track_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_18_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_19_ccff_tail),
		.mem_out(mem_out[158:159]),
		.mem_outb(mem_outb[158:159]));

	sb_mux_size2_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_19_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_20_ccff_tail),
		.mem_out(mem_out[160:161]),
		.mem_outb(mem_outb[160:161]));

	sb_mux_size2_mem mem_bottom_track_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_20_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_21_ccff_tail),
		.mem_out(mem_out[162:163]),
		.mem_outb(mem_outb[162:163]));

	sb_mux_size2_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_21_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_22_ccff_tail),
		.mem_out(mem_out[164:165]),
		.mem_outb(mem_outb[164:165]));

	sb_mux_size2_mem mem_bottom_track_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_22_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_23_ccff_tail),
		.mem_out(mem_out[166:167]),
		.mem_outb(mem_outb[166:167]));

	sb_mux_size2_mem mem_bottom_track_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_23_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_24_ccff_tail),
		.mem_out(mem_out[168:169]),
		.mem_outb(mem_outb[168:169]));

	sb_mux_size2_mem mem_bottom_track_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_24_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_25_ccff_tail),
		.mem_out(mem_out[170:171]),
		.mem_outb(mem_outb[170:171]));

	sb_mux_size2_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_25_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_26_ccff_tail),
		.mem_out(mem_out[172:173]),
		.mem_outb(mem_outb[172:173]));

	sb_mux_size2_mem mem_bottom_track_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_26_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_27_ccff_tail),
		.mem_out(mem_out[174:175]),
		.mem_outb(mem_outb[174:175]));

	sb_mux_size2_mem mem_bottom_track_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_27_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_28_ccff_tail),
		.mem_out(mem_out[176:177]),
		.mem_outb(mem_outb[176:177]));

	sb_mux_size2_mem mem_bottom_track_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_28_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_29_ccff_tail),
		.mem_out(mem_out[178:179]),
		.mem_outb(mem_outb[178:179]));

endmodule
// ----- END Verilog module for sb_4__config_group_mem_size244 -----




// ----- Verilog module for sb_6__config_group_mem_size340 -----
module sb_6__config_group_mem_size340(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:339] mem_out;
//----- OUTPUT PORTS -----
output [0:339] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size10_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size10_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size10_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size10_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_3_ccff_tail),
		.mem_out(mem_out[22:25]),
		.mem_outb(mem_outb[22:25]));

	sb_mux_size10_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_4_ccff_tail),
		.mem_out(mem_out[26:29]),
		.mem_outb(mem_outb[26:29]));

	sb_mux_size10_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_5_ccff_tail),
		.mem_out(mem_out[30:33]),
		.mem_outb(mem_outb[30:33]));

	sb_mux_size10_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_6_ccff_tail),
		.mem_out(mem_out[170:173]),
		.mem_outb(mem_outb[170:173]));

	sb_mux_size10_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_7_ccff_tail),
		.mem_out(mem_out[174:177]),
		.mem_outb(mem_outb[174:177]));

	sb_mux_size10_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_8_ccff_tail),
		.mem_out(mem_out[178:181]),
		.mem_outb(mem_outb[178:181]));

	sb_mux_size10_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_9_ccff_tail),
		.mem_out(mem_out[192:195]),
		.mem_outb(mem_outb[192:195]));

	sb_mux_size10_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_10_ccff_tail),
		.mem_out(mem_out[196:199]),
		.mem_outb(mem_outb[196:199]));

	sb_mux_size10_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_11_ccff_tail),
		.mem_out(mem_out[200:203]),
		.mem_outb(mem_outb[200:203]));

	sb_mux_size9_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size9_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[126:129]),
		.mem_outb(mem_outb[126:129]));

	sb_mux_size9_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_2_ccff_tail),
		.mem_out(mem_out[130:133]),
		.mem_outb(mem_outb[130:133]));

	sb_mux_size9_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_3_ccff_tail),
		.mem_out(mem_out[148:151]),
		.mem_outb(mem_outb[148:151]));

	sb_mux_size9_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_4_ccff_tail),
		.mem_out(mem_out[152:155]),
		.mem_outb(mem_outb[152:155]));

	sb_mux_size9_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_5_ccff_tail),
		.mem_out(mem_out[156:159]),
		.mem_outb(mem_outb[156:159]));

	sb_mux_size9_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_6_ccff_tail),
		.mem_out(mem_out[160:163]),
		.mem_outb(mem_outb[160:163]));

	sb_mux_size9_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_7_ccff_tail),
		.mem_out(mem_out[182:185]),
		.mem_outb(mem_outb[182:185]));

	sb_mux_size9_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_8_ccff_tail),
		.mem_out(mem_out[296:299]),
		.mem_outb(mem_outb[296:299]));

	sb_mux_size9_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_9_ccff_tail),
		.mem_out(mem_out[300:303]),
		.mem_outb(mem_outb[300:303]));

	sb_mux_size9_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_10_ccff_tail),
		.mem_out(mem_out[318:321]),
		.mem_outb(mem_outb[318:321]));

	sb_mux_size9_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_11_ccff_tail),
		.mem_out(mem_out[322:325]),
		.mem_outb(mem_outb[322:325]));

	sb_mux_size9_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_12_ccff_tail),
		.mem_out(mem_out[326:329]),
		.mem_outb(mem_outb[326:329]));

	sb_mux_size9_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_13_ccff_tail),
		.mem_out(mem_out[330:333]),
		.mem_outb(mem_outb[330:333]));

	sb_mux_size7_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_0_ccff_tail),
		.mem_out(mem_out[16:18]),
		.mem_outb(mem_outb[16:18]));

	sb_mux_size7_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_1_ccff_tail),
		.mem_out(mem_out[19:21]),
		.mem_outb(mem_outb[19:21]));

	sb_mux_size7_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_2_ccff_tail),
		.mem_out(mem_out[134:136]),
		.mem_outb(mem_outb[134:136]));

	sb_mux_size7_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_3_ccff_tail),
		.mem_out(mem_out[137:139]),
		.mem_outb(mem_outb[137:139]));

	sb_mux_size7_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_4_ccff_tail),
		.mem_out(mem_out[164:166]),
		.mem_outb(mem_outb[164:166]));

	sb_mux_size7_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_5_ccff_tail),
		.mem_out(mem_out[167:169]),
		.mem_outb(mem_outb[167:169]));

	sb_mux_size7_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_6_ccff_tail),
		.mem_out(mem_out[186:188]),
		.mem_outb(mem_outb[186:188]));

	sb_mux_size7_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_7_ccff_tail),
		.mem_out(mem_out[189:191]),
		.mem_outb(mem_outb[189:191]));

	sb_mux_size7_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_8_ccff_tail),
		.mem_out(mem_out[304:306]),
		.mem_outb(mem_outb[304:306]));

	sb_mux_size7_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_9_ccff_tail),
		.mem_out(mem_out[307:309]),
		.mem_outb(mem_outb[307:309]));

	sb_mux_size7_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_10_ccff_tail),
		.mem_out(mem_out[334:336]),
		.mem_outb(mem_outb[334:336]));

	sb_mux_size7_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_10_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[337:339]),
		.mem_outb(mem_outb[337:339]));

	sb_mux_size8_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[34:37]),
		.mem_outb(mem_outb[34:37]));

	sb_mux_size8_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[38:41]),
		.mem_outb(mem_outb[38:41]));

	sb_mux_size8_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[42:45]),
		.mem_outb(mem_outb[42:45]));

	sb_mux_size8_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[46:49]),
		.mem_outb(mem_outb[46:49]));

	sb_mux_size8_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[50:53]),
		.mem_outb(mem_outb[50:53]));

	sb_mux_size8_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[204:207]),
		.mem_outb(mem_outb[204:207]));

	sb_mux_size8_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[208:211]),
		.mem_outb(mem_outb[208:211]));

	sb_mux_size8_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[212:215]),
		.mem_outb(mem_outb[212:215]));

	sb_mux_size8_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[216:219]),
		.mem_outb(mem_outb[216:219]));

	sb_mux_size8_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[220:223]),
		.mem_outb(mem_outb[220:223]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[54:55]),
		.mem_outb(mem_outb[54:55]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[64:65]),
		.mem_outb(mem_outb[64:65]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[66:67]),
		.mem_outb(mem_outb[66:67]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[68:69]),
		.mem_outb(mem_outb[68:69]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[70:71]),
		.mem_outb(mem_outb[70:71]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[72:73]),
		.mem_outb(mem_outb[72:73]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[74:75]),
		.mem_outb(mem_outb[74:75]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[76:77]),
		.mem_outb(mem_outb[76:77]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[78:79]),
		.mem_outb(mem_outb[78:79]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[80:81]),
		.mem_outb(mem_outb[80:81]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[82:83]),
		.mem_outb(mem_outb[82:83]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[84:85]),
		.mem_outb(mem_outb[84:85]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[86:87]),
		.mem_outb(mem_outb[86:87]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[88:89]),
		.mem_outb(mem_outb[88:89]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[94:95]),
		.mem_outb(mem_outb[94:95]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[96:97]),
		.mem_outb(mem_outb[96:97]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[98:99]),
		.mem_outb(mem_outb[98:99]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[116:117]),
		.mem_outb(mem_outb[116:117]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[224:225]),
		.mem_outb(mem_outb[224:225]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[226:227]),
		.mem_outb(mem_outb[226:227]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[228:229]),
		.mem_outb(mem_outb[228:229]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[230:231]),
		.mem_outb(mem_outb[230:231]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[232:233]),
		.mem_outb(mem_outb[232:233]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[234:235]),
		.mem_outb(mem_outb[234:235]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[236:237]),
		.mem_outb(mem_outb[236:237]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[238:239]),
		.mem_outb(mem_outb[238:239]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[240:241]),
		.mem_outb(mem_outb[240:241]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[242:243]),
		.mem_outb(mem_outb[242:243]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[244:245]),
		.mem_outb(mem_outb[244:245]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[246:247]),
		.mem_outb(mem_outb[246:247]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[248:249]),
		.mem_outb(mem_outb[248:249]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[250:251]),
		.mem_outb(mem_outb[250:251]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[252:253]),
		.mem_outb(mem_outb[252:253]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[254:255]),
		.mem_outb(mem_outb[254:255]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[256:257]),
		.mem_outb(mem_outb[256:257]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[258:259]),
		.mem_outb(mem_outb[258:259]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[260:261]),
		.mem_outb(mem_outb[260:261]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[262:263]),
		.mem_outb(mem_outb[262:263]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[264:265]),
		.mem_outb(mem_outb[264:265]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[266:267]),
		.mem_outb(mem_outb[266:267]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[268:269]),
		.mem_outb(mem_outb[268:269]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[270:271]),
		.mem_outb(mem_outb[270:271]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[272:273]),
		.mem_outb(mem_outb[272:273]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[274:275]),
		.mem_outb(mem_outb[274:275]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[276:277]),
		.mem_outb(mem_outb[276:277]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[278:279]),
		.mem_outb(mem_outb[278:279]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[280:281]),
		.mem_outb(mem_outb[280:281]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[282:283]),
		.mem_outb(mem_outb[282:283]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[284:285]),
		.mem_outb(mem_outb[284:285]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[286:287]),
		.mem_outb(mem_outb[286:287]));

	sb_mux_size11_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[118:121]),
		.mem_outb(mem_outb[118:121]));

	sb_mux_size11_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[122:125]),
		.mem_outb(mem_outb[122:125]));

	sb_mux_size11_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[140:143]),
		.mem_outb(mem_outb[140:143]));

	sb_mux_size11_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[144:147]),
		.mem_outb(mem_outb[144:147]));

	sb_mux_size11_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_4_ccff_tail),
		.mem_out(mem_out[288:291]),
		.mem_outb(mem_outb[288:291]));

	sb_mux_size11_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_5_ccff_tail),
		.mem_out(mem_out[292:295]),
		.mem_outb(mem_outb[292:295]));

	sb_mux_size11_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_6_ccff_tail),
		.mem_out(mem_out[310:313]),
		.mem_outb(mem_outb[310:313]));

	sb_mux_size11_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_7_ccff_tail),
		.mem_out(mem_out[314:317]),
		.mem_outb(mem_outb[314:317]));

endmodule
// ----- END Verilog module for sb_6__config_group_mem_size340 -----




// ----- Verilog module for sb_7__config_group_mem_size358 -----
module sb_7__config_group_mem_size358(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:357] mem_out;
//----- OUTPUT PORTS -----
output [0:357] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size13_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size13_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size13_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size13_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size13_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_3_ccff_tail),
		.mem_out(mem_out[120:123]),
		.mem_outb(mem_outb[120:123]));

	sb_mux_size13_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_4_ccff_tail),
		.mem_out(mem_out[124:127]),
		.mem_outb(mem_outb[124:127]));

	sb_mux_size13_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_5_ccff_tail),
		.mem_out(mem_out[128:131]),
		.mem_outb(mem_outb[128:131]));

	sb_mux_size13_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_6_ccff_tail),
		.mem_out(mem_out[132:135]),
		.mem_outb(mem_outb[132:135]));

	sb_mux_size13_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_7_ccff_tail),
		.mem_out(mem_out[159:162]),
		.mem_outb(mem_outb[159:162]));

	sb_mux_size13_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_8_ccff_tail),
		.mem_out(mem_out[163:166]),
		.mem_outb(mem_outb[163:166]));

	sb_mux_size13_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_9_ccff_tail),
		.mem_out(mem_out[167:170]),
		.mem_outb(mem_outb[167:170]));

	sb_mux_size13_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_10_ccff_tail),
		.mem_out(mem_out[179:182]),
		.mem_outb(mem_outb[179:182]));

	sb_mux_size13_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_11_ccff_tail),
		.mem_out(mem_out[183:186]),
		.mem_outb(mem_outb[183:186]));

	sb_mux_size13_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_12_ccff_tail),
		.mem_out(mem_out[187:190]),
		.mem_outb(mem_outb[187:190]));

	sb_mux_size13_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_13_ccff_tail),
		.mem_out(mem_out[299:302]),
		.mem_outb(mem_outb[299:302]));

	sb_mux_size13_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_14_ccff_tail),
		.mem_out(mem_out[303:306]),
		.mem_outb(mem_outb[303:306]));

	sb_mux_size13_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_15_ccff_tail),
		.mem_out(mem_out[307:310]),
		.mem_outb(mem_outb[307:310]));

	sb_mux_size13_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_15_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_16_ccff_tail),
		.mem_out(mem_out[311:314]),
		.mem_outb(mem_outb[311:314]));

	sb_mux_size13_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_17_ccff_tail),
		.mem_out(mem_out[338:341]),
		.mem_outb(mem_outb[338:341]));

	sb_mux_size13_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_17_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_18_ccff_tail),
		.mem_out(mem_out[342:345]),
		.mem_outb(mem_outb[342:345]));

	sb_mux_size13_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_18_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_19_ccff_tail),
		.mem_out(mem_out[346:349]),
		.mem_outb(mem_outb[346:349]));

	sb_mux_size11_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size11_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[36:39]),
		.mem_outb(mem_outb[36:39]));

	sb_mux_size11_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[40:43]),
		.mem_outb(mem_outb[40:43]));

	sb_mux_size11_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[44:47]),
		.mem_outb(mem_outb[44:47]));

	sb_mux_size11_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_4_ccff_tail),
		.mem_out(mem_out[48:51]),
		.mem_outb(mem_outb[48:51]));

	sb_mux_size11_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_5_ccff_tail),
		.mem_out(mem_out[52:55]),
		.mem_outb(mem_outb[52:55]));

	sb_mux_size11_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_6_ccff_tail),
		.mem_out(mem_out[136:139]),
		.mem_outb(mem_outb[136:139]));

	sb_mux_size11_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_7_ccff_tail),
		.mem_out(mem_out[140:143]),
		.mem_outb(mem_outb[140:143]));

	sb_mux_size11_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_8_ccff_tail),
		.mem_out(mem_out[171:174]),
		.mem_outb(mem_outb[171:174]));

	sb_mux_size11_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_9_ccff_tail),
		.mem_out(mem_out[175:178]),
		.mem_outb(mem_outb[175:178]));

	sb_mux_size11_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_10_ccff_tail),
		.mem_out(mem_out[191:194]),
		.mem_outb(mem_outb[191:194]));

	sb_mux_size11_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_11_ccff_tail),
		.mem_out(mem_out[215:218]),
		.mem_outb(mem_outb[215:218]));

	sb_mux_size11_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_12_ccff_tail),
		.mem_out(mem_out[219:222]),
		.mem_outb(mem_outb[219:222]));

	sb_mux_size11_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_13_ccff_tail),
		.mem_out(mem_out[223:226]),
		.mem_outb(mem_outb[223:226]));

	sb_mux_size11_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_14_ccff_tail),
		.mem_out(mem_out[227:230]),
		.mem_outb(mem_outb[227:230]));

	sb_mux_size11_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_15_ccff_tail),
		.mem_out(mem_out[231:234]),
		.mem_outb(mem_outb[231:234]));

	sb_mux_size11_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_16_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_16_ccff_tail),
		.mem_out(mem_out[315:318]),
		.mem_outb(mem_outb[315:318]));

	sb_mux_size11_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_16_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_17_ccff_tail),
		.mem_out(mem_out[319:322]),
		.mem_outb(mem_outb[319:322]));

	sb_mux_size11_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_19_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_18_ccff_tail),
		.mem_out(mem_out[350:353]),
		.mem_outb(mem_outb[350:353]));

	sb_mux_size11_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_18_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[354:357]),
		.mem_outb(mem_outb[354:357]));

	sb_mux_size9_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[16:19]),
		.mem_outb(mem_outb[16:19]));

	sb_mux_size9_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[20:23]),
		.mem_outb(mem_outb[20:23]));

	sb_mux_size9_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_2_ccff_tail),
		.mem_out(mem_out[195:198]),
		.mem_outb(mem_outb[195:198]));

	sb_mux_size9_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_3_ccff_tail),
		.mem_out(mem_out[199:202]),
		.mem_outb(mem_outb[199:202]));

	sb_mux_size15_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_0_ccff_tail),
		.mem_out(mem_out[24:27]),
		.mem_outb(mem_outb[24:27]));

	sb_mux_size15_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_1_ccff_tail),
		.mem_out(mem_out[28:31]),
		.mem_outb(mem_outb[28:31]));

	sb_mux_size15_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_2_ccff_tail),
		.mem_out(mem_out[32:35]),
		.mem_outb(mem_outb[32:35]));

	sb_mux_size15_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_3_ccff_tail),
		.mem_out(mem_out[203:206]),
		.mem_outb(mem_outb[203:206]));

	sb_mux_size15_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_4_ccff_tail),
		.mem_out(mem_out[207:210]),
		.mem_outb(mem_outb[207:210]));

	sb_mux_size15_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_5_ccff_tail),
		.mem_out(mem_out[211:214]),
		.mem_outb(mem_outb[211:214]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[64:65]),
		.mem_outb(mem_outb[64:65]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[66:67]),
		.mem_outb(mem_outb[66:67]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[68:69]),
		.mem_outb(mem_outb[68:69]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[70:71]),
		.mem_outb(mem_outb[70:71]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[72:73]),
		.mem_outb(mem_outb[72:73]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[74:75]),
		.mem_outb(mem_outb[74:75]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[76:77]),
		.mem_outb(mem_outb[76:77]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[78:79]),
		.mem_outb(mem_outb[78:79]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[80:81]),
		.mem_outb(mem_outb[80:81]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[82:83]),
		.mem_outb(mem_outb[82:83]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[84:85]),
		.mem_outb(mem_outb[84:85]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[86:87]),
		.mem_outb(mem_outb[86:87]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[88:89]),
		.mem_outb(mem_outb[88:89]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[94:95]),
		.mem_outb(mem_outb[94:95]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[96:97]),
		.mem_outb(mem_outb[96:97]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[98:99]),
		.mem_outb(mem_outb[98:99]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[116:117]),
		.mem_outb(mem_outb[116:117]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[118:119]),
		.mem_outb(mem_outb[118:119]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[235:236]),
		.mem_outb(mem_outb[235:236]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[237:238]),
		.mem_outb(mem_outb[237:238]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[239:240]),
		.mem_outb(mem_outb[239:240]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[241:242]),
		.mem_outb(mem_outb[241:242]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[243:244]),
		.mem_outb(mem_outb[243:244]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[245:246]),
		.mem_outb(mem_outb[245:246]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[247:248]),
		.mem_outb(mem_outb[247:248]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[249:250]),
		.mem_outb(mem_outb[249:250]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[251:252]),
		.mem_outb(mem_outb[251:252]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[253:254]),
		.mem_outb(mem_outb[253:254]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[255:256]),
		.mem_outb(mem_outb[255:256]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[257:258]),
		.mem_outb(mem_outb[257:258]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[259:260]),
		.mem_outb(mem_outb[259:260]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[261:262]),
		.mem_outb(mem_outb[261:262]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[263:264]),
		.mem_outb(mem_outb[263:264]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[265:266]),
		.mem_outb(mem_outb[265:266]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[267:268]),
		.mem_outb(mem_outb[267:268]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[269:270]),
		.mem_outb(mem_outb[269:270]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[271:272]),
		.mem_outb(mem_outb[271:272]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[273:274]),
		.mem_outb(mem_outb[273:274]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[275:276]),
		.mem_outb(mem_outb[275:276]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[277:278]),
		.mem_outb(mem_outb[277:278]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[279:280]),
		.mem_outb(mem_outb[279:280]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[281:282]),
		.mem_outb(mem_outb[281:282]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[283:284]),
		.mem_outb(mem_outb[283:284]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[285:286]),
		.mem_outb(mem_outb[285:286]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[287:288]),
		.mem_outb(mem_outb[287:288]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[289:290]),
		.mem_outb(mem_outb[289:290]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[291:292]),
		.mem_outb(mem_outb[291:292]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[293:294]),
		.mem_outb(mem_outb[293:294]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[295:296]),
		.mem_outb(mem_outb[295:296]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[297:298]),
		.mem_outb(mem_outb[297:298]));

	sb_mux_size17_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_0_ccff_tail),
		.mem_out(mem_out[144:148]),
		.mem_outb(mem_outb[144:148]));

	sb_mux_size17_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_1_ccff_tail),
		.mem_out(mem_out[149:153]),
		.mem_outb(mem_outb[149:153]));

	sb_mux_size17_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_2_ccff_tail),
		.mem_out(mem_out[154:158]),
		.mem_outb(mem_outb[154:158]));

	sb_mux_size17_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_17_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_3_ccff_tail),
		.mem_out(mem_out[323:327]),
		.mem_outb(mem_outb[323:327]));

	sb_mux_size17_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_4_ccff_tail),
		.mem_out(mem_out[328:332]),
		.mem_outb(mem_outb[328:332]));

	sb_mux_size17_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_5_ccff_tail),
		.mem_out(mem_out[333:337]),
		.mem_outb(mem_outb[333:337]));

endmodule
// ----- END Verilog module for sb_7__config_group_mem_size358 -----




// ----- Verilog module for sb_8__config_group_mem_size360 -----
module sb_8__config_group_mem_size360(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:359] mem_out;
//----- OUTPUT PORTS -----
output [0:359] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size10_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size10_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size10_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size10_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_3_ccff_tail),
		.mem_out(mem_out[22:25]),
		.mem_outb(mem_outb[22:25]));

	sb_mux_size10_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_4_ccff_tail),
		.mem_out(mem_out[26:29]),
		.mem_outb(mem_outb[26:29]));

	sb_mux_size10_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_5_ccff_tail),
		.mem_out(mem_out[30:33]),
		.mem_outb(mem_outb[30:33]));

	sb_mux_size10_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_6_ccff_tail),
		.mem_out(mem_out[180:183]),
		.mem_outb(mem_outb[180:183]));

	sb_mux_size10_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_7_ccff_tail),
		.mem_out(mem_out[184:187]),
		.mem_outb(mem_outb[184:187]));

	sb_mux_size10_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_8_ccff_tail),
		.mem_out(mem_out[188:191]),
		.mem_outb(mem_outb[188:191]));

	sb_mux_size10_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_9_ccff_tail),
		.mem_out(mem_out[202:205]),
		.mem_outb(mem_outb[202:205]));

	sb_mux_size10_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_10_ccff_tail),
		.mem_out(mem_out[206:209]),
		.mem_outb(mem_outb[206:209]));

	sb_mux_size10_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_11_ccff_tail),
		.mem_out(mem_out[210:213]),
		.mem_outb(mem_outb[210:213]));

	sb_mux_size9_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size9_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[192:195]),
		.mem_outb(mem_outb[192:195]));

	sb_mux_size7_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_0_ccff_tail),
		.mem_out(mem_out[16:18]),
		.mem_outb(mem_outb[16:18]));

	sb_mux_size7_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_1_ccff_tail),
		.mem_out(mem_out[19:21]),
		.mem_outb(mem_outb[19:21]));

	sb_mux_size7_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_2_ccff_tail),
		.mem_out(mem_out[196:198]),
		.mem_outb(mem_outb[196:198]));

	sb_mux_size7_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_3_ccff_tail),
		.mem_out(mem_out[199:201]),
		.mem_outb(mem_outb[199:201]));

	sb_mux_size8_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[34:37]),
		.mem_outb(mem_outb[34:37]));

	sb_mux_size8_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[38:41]),
		.mem_outb(mem_outb[38:41]));

	sb_mux_size8_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[42:45]),
		.mem_outb(mem_outb[42:45]));

	sb_mux_size8_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[46:49]),
		.mem_outb(mem_outb[46:49]));

	sb_mux_size8_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[50:53]),
		.mem_outb(mem_outb[50:53]));

	sb_mux_size8_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[214:217]),
		.mem_outb(mem_outb[214:217]));

	sb_mux_size8_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[218:221]),
		.mem_outb(mem_outb[218:221]));

	sb_mux_size8_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[222:225]),
		.mem_outb(mem_outb[222:225]));

	sb_mux_size8_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[226:229]),
		.mem_outb(mem_outb[226:229]));

	sb_mux_size8_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[230:233]),
		.mem_outb(mem_outb[230:233]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[54:55]),
		.mem_outb(mem_outb[54:55]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[64:65]),
		.mem_outb(mem_outb[64:65]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[66:67]),
		.mem_outb(mem_outb[66:67]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[68:69]),
		.mem_outb(mem_outb[68:69]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[70:71]),
		.mem_outb(mem_outb[70:71]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[72:73]),
		.mem_outb(mem_outb[72:73]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[74:75]),
		.mem_outb(mem_outb[74:75]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[76:77]),
		.mem_outb(mem_outb[76:77]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[78:79]),
		.mem_outb(mem_outb[78:79]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[80:81]),
		.mem_outb(mem_outb[80:81]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[82:83]),
		.mem_outb(mem_outb[82:83]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[84:85]),
		.mem_outb(mem_outb[84:85]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[86:87]),
		.mem_outb(mem_outb[86:87]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[88:89]),
		.mem_outb(mem_outb[88:89]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[94:95]),
		.mem_outb(mem_outb[94:95]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[96:97]),
		.mem_outb(mem_outb[96:97]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[98:99]),
		.mem_outb(mem_outb[98:99]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[116:117]),
		.mem_outb(mem_outb[116:117]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[234:235]),
		.mem_outb(mem_outb[234:235]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[236:237]),
		.mem_outb(mem_outb[236:237]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[238:239]),
		.mem_outb(mem_outb[238:239]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[240:241]),
		.mem_outb(mem_outb[240:241]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[242:243]),
		.mem_outb(mem_outb[242:243]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[244:245]),
		.mem_outb(mem_outb[244:245]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[246:247]),
		.mem_outb(mem_outb[246:247]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[248:249]),
		.mem_outb(mem_outb[248:249]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[250:251]),
		.mem_outb(mem_outb[250:251]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[252:253]),
		.mem_outb(mem_outb[252:253]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[254:255]),
		.mem_outb(mem_outb[254:255]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[256:257]),
		.mem_outb(mem_outb[256:257]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[258:259]),
		.mem_outb(mem_outb[258:259]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[260:261]),
		.mem_outb(mem_outb[260:261]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[262:263]),
		.mem_outb(mem_outb[262:263]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[264:265]),
		.mem_outb(mem_outb[264:265]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[266:267]),
		.mem_outb(mem_outb[266:267]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[268:269]),
		.mem_outb(mem_outb[268:269]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[270:271]),
		.mem_outb(mem_outb[270:271]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[272:273]),
		.mem_outb(mem_outb[272:273]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[274:275]),
		.mem_outb(mem_outb[274:275]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[276:277]),
		.mem_outb(mem_outb[276:277]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[278:279]),
		.mem_outb(mem_outb[278:279]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[280:281]),
		.mem_outb(mem_outb[280:281]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[282:283]),
		.mem_outb(mem_outb[282:283]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[284:285]),
		.mem_outb(mem_outb[284:285]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[286:287]),
		.mem_outb(mem_outb[286:287]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[288:289]),
		.mem_outb(mem_outb[288:289]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[290:291]),
		.mem_outb(mem_outb[290:291]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[292:293]),
		.mem_outb(mem_outb[292:293]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[294:295]),
		.mem_outb(mem_outb[294:295]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[296:297]),
		.mem_outb(mem_outb[296:297]));

	sb_mux_size17_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_0_ccff_tail),
		.mem_out(mem_out[118:122]),
		.mem_outb(mem_outb[118:122]));

	sb_mux_size17_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_1_ccff_tail),
		.mem_out(mem_out[123:127]),
		.mem_outb(mem_outb[123:127]));

	sb_mux_size17_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size21_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_2_ccff_tail),
		.mem_out(mem_out[159:163]),
		.mem_outb(mem_outb[159:163]));

	sb_mux_size17_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_3_ccff_tail),
		.mem_out(mem_out[298:302]),
		.mem_outb(mem_outb[298:302]));

	sb_mux_size17_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_4_ccff_tail),
		.mem_out(mem_out[303:307]),
		.mem_outb(mem_outb[303:307]));

	sb_mux_size17_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size21_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size17_mem_5_ccff_tail),
		.mem_out(mem_out[339:343]),
		.mem_outb(mem_outb[339:343]));

	sb_mux_size15_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_0_ccff_tail),
		.mem_out(mem_out[128:131]),
		.mem_outb(mem_outb[128:131]));

	sb_mux_size15_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_1_ccff_tail),
		.mem_out(mem_out[132:135]),
		.mem_outb(mem_outb[132:135]));

	sb_mux_size15_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_2_ccff_tail),
		.mem_out(mem_out[164:167]),
		.mem_outb(mem_outb[164:167]));

	sb_mux_size15_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_3_ccff_tail),
		.mem_out(mem_out[168:171]),
		.mem_outb(mem_outb[168:171]));

	sb_mux_size15_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_4_ccff_tail),
		.mem_out(mem_out[172:175]),
		.mem_outb(mem_outb[172:175]));

	sb_mux_size15_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_5_ccff_tail),
		.mem_out(mem_out[176:179]),
		.mem_outb(mem_outb[176:179]));

	sb_mux_size15_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_6_ccff_tail),
		.mem_out(mem_out[308:311]),
		.mem_outb(mem_outb[308:311]));

	sb_mux_size15_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_7_ccff_tail),
		.mem_out(mem_out[312:315]),
		.mem_outb(mem_outb[312:315]));

	sb_mux_size15_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size17_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_8_ccff_tail),
		.mem_out(mem_out[344:347]),
		.mem_outb(mem_outb[344:347]));

	sb_mux_size15_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_9_ccff_tail),
		.mem_out(mem_out[348:351]),
		.mem_outb(mem_outb[348:351]));

	sb_mux_size15_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_10_ccff_tail),
		.mem_out(mem_out[352:355]),
		.mem_outb(mem_outb[352:355]));

	sb_mux_size15_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_10_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[356:359]),
		.mem_outb(mem_outb[356:359]));

	sb_mux_size13_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_0_ccff_tail),
		.mem_out(mem_out[136:139]),
		.mem_outb(mem_outb[136:139]));

	sb_mux_size13_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_1_ccff_tail),
		.mem_out(mem_out[140:143]),
		.mem_outb(mem_outb[140:143]));

	sb_mux_size13_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_2_ccff_tail),
		.mem_out(mem_out[316:319]),
		.mem_outb(mem_outb[316:319]));

	sb_mux_size13_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_3_ccff_tail),
		.mem_out(mem_out[320:323]),
		.mem_outb(mem_outb[320:323]));

	sb_mux_size23_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size23_mem_0_ccff_tail),
		.mem_out(mem_out[144:148]),
		.mem_outb(mem_outb[144:148]));

	sb_mux_size23_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size23_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size23_mem_1_ccff_tail),
		.mem_out(mem_out[149:153]),
		.mem_outb(mem_outb[149:153]));

	sb_mux_size23_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size23_mem_2_ccff_tail),
		.mem_out(mem_out[324:328]),
		.mem_outb(mem_outb[324:328]));

	sb_mux_size23_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size23_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size23_mem_3_ccff_tail),
		.mem_out(mem_out[329:333]),
		.mem_outb(mem_outb[329:333]));

	sb_mux_size21_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size23_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size21_mem_0_ccff_tail),
		.mem_out(mem_out[154:158]),
		.mem_outb(mem_outb[154:158]));

	sb_mux_size21_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size23_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size21_mem_1_ccff_tail),
		.mem_out(mem_out[334:338]),
		.mem_outb(mem_outb[334:338]));

endmodule
// ----- END Verilog module for sb_8__config_group_mem_size360 -----




// ----- Verilog module for sb_10__config_group_mem_size336 -----
module sb_10__config_group_mem_size336(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:335] mem_out;
//----- OUTPUT PORTS -----
output [0:335] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size11_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size11_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size11_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size11_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size11_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_4_ccff_tail),
		.mem_out(mem_out[168:171]),
		.mem_outb(mem_outb[168:171]));

	sb_mux_size11_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_5_ccff_tail),
		.mem_out(mem_out[172:175]),
		.mem_outb(mem_outb[172:175]));

	sb_mux_size11_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_6_ccff_tail),
		.mem_out(mem_out[176:179]),
		.mem_outb(mem_outb[176:179]));

	sb_mux_size11_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_7_ccff_tail),
		.mem_out(mem_out[180:183]),
		.mem_outb(mem_outb[180:183]));

	sb_mux_size9_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[16:19]),
		.mem_outb(mem_outb[16:19]));

	sb_mux_size9_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[48:51]),
		.mem_outb(mem_outb[48:51]));

	sb_mux_size9_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_2_ccff_tail),
		.mem_out(mem_out[52:55]),
		.mem_outb(mem_outb[52:55]));

	sb_mux_size9_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_3_ccff_tail),
		.mem_out(mem_out[120:123]),
		.mem_outb(mem_outb[120:123]));

	sb_mux_size9_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_4_ccff_tail),
		.mem_out(mem_out[124:127]),
		.mem_outb(mem_outb[124:127]));

	sb_mux_size9_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_5_ccff_tail),
		.mem_out(mem_out[184:187]),
		.mem_outb(mem_outb[184:187]));

	sb_mux_size9_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_6_ccff_tail),
		.mem_out(mem_out[216:219]),
		.mem_outb(mem_outb[216:219]));

	sb_mux_size9_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_7_ccff_tail),
		.mem_out(mem_out[220:223]),
		.mem_outb(mem_outb[220:223]));

	sb_mux_size9_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_8_ccff_tail),
		.mem_out(mem_out[288:291]),
		.mem_outb(mem_outb[288:291]));

	sb_mux_size9_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_9_ccff_tail),
		.mem_out(mem_out[292:295]),
		.mem_outb(mem_outb[292:295]));

	sb_mux_size8_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[20:23]),
		.mem_outb(mem_outb[20:23]));

	sb_mux_size8_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[128:131]),
		.mem_outb(mem_outb[128:131]));

	sb_mux_size8_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[132:135]),
		.mem_outb(mem_outb[132:135]));

	sb_mux_size8_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[142:145]),
		.mem_outb(mem_outb[142:145]));

	sb_mux_size8_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[146:149]),
		.mem_outb(mem_outb[146:149]));

	sb_mux_size8_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[188:191]),
		.mem_outb(mem_outb[188:191]));

	sb_mux_size8_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[296:299]),
		.mem_outb(mem_outb[296:299]));

	sb_mux_size8_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[300:303]),
		.mem_outb(mem_outb[300:303]));

	sb_mux_size8_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[310:313]),
		.mem_outb(mem_outb[310:313]));

	sb_mux_size8_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[314:317]),
		.mem_outb(mem_outb[314:317]));

	sb_mux_size13_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_0_ccff_tail),
		.mem_out(mem_out[24:27]),
		.mem_outb(mem_outb[24:27]));

	sb_mux_size13_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_1_ccff_tail),
		.mem_out(mem_out[28:31]),
		.mem_outb(mem_outb[28:31]));

	sb_mux_size13_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_2_ccff_tail),
		.mem_out(mem_out[192:195]),
		.mem_outb(mem_outb[192:195]));

	sb_mux_size13_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_3_ccff_tail),
		.mem_out(mem_out[196:199]),
		.mem_outb(mem_outb[196:199]));

	sb_mux_size12_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size12_mem_0_ccff_tail),
		.mem_out(mem_out[32:35]),
		.mem_outb(mem_outb[32:35]));

	sb_mux_size12_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size12_mem_1_ccff_tail),
		.mem_out(mem_out[200:203]),
		.mem_outb(mem_outb[200:203]));

	sb_mux_size10_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size12_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[36:39]),
		.mem_outb(mem_outb[36:39]));

	sb_mux_size10_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[40:43]),
		.mem_outb(mem_outb[40:43]));

	sb_mux_size10_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_2_ccff_tail),
		.mem_out(mem_out[44:47]),
		.mem_outb(mem_outb[44:47]));

	sb_mux_size10_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size12_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_3_ccff_tail),
		.mem_out(mem_out[204:207]),
		.mem_outb(mem_outb[204:207]));

	sb_mux_size10_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_4_ccff_tail),
		.mem_out(mem_out[208:211]),
		.mem_outb(mem_outb[208:211]));

	sb_mux_size10_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_5_ccff_tail),
		.mem_out(mem_out[212:215]),
		.mem_outb(mem_outb[212:215]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[56:57]),
		.mem_outb(mem_outb[56:57]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[58:59]),
		.mem_outb(mem_outb[58:59]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[60:61]),
		.mem_outb(mem_outb[60:61]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[62:63]),
		.mem_outb(mem_outb[62:63]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[64:65]),
		.mem_outb(mem_outb[64:65]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[66:67]),
		.mem_outb(mem_outb[66:67]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[68:69]),
		.mem_outb(mem_outb[68:69]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[70:71]),
		.mem_outb(mem_outb[70:71]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[72:73]),
		.mem_outb(mem_outb[72:73]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[74:75]),
		.mem_outb(mem_outb[74:75]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[76:77]),
		.mem_outb(mem_outb[76:77]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[78:79]),
		.mem_outb(mem_outb[78:79]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[80:81]),
		.mem_outb(mem_outb[80:81]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[82:83]),
		.mem_outb(mem_outb[82:83]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[84:85]),
		.mem_outb(mem_outb[84:85]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[86:87]),
		.mem_outb(mem_outb[86:87]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[88:89]),
		.mem_outb(mem_outb[88:89]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[90:91]),
		.mem_outb(mem_outb[90:91]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[92:93]),
		.mem_outb(mem_outb[92:93]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[94:95]),
		.mem_outb(mem_outb[94:95]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[96:97]),
		.mem_outb(mem_outb[96:97]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[98:99]),
		.mem_outb(mem_outb[98:99]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[100:101]),
		.mem_outb(mem_outb[100:101]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[102:103]),
		.mem_outb(mem_outb[102:103]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[104:105]),
		.mem_outb(mem_outb[104:105]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[106:107]),
		.mem_outb(mem_outb[106:107]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[108:109]),
		.mem_outb(mem_outb[108:109]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[110:111]),
		.mem_outb(mem_outb[110:111]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[112:113]),
		.mem_outb(mem_outb[112:113]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[114:115]),
		.mem_outb(mem_outb[114:115]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[116:117]),
		.mem_outb(mem_outb[116:117]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[118:119]),
		.mem_outb(mem_outb[118:119]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[224:225]),
		.mem_outb(mem_outb[224:225]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[226:227]),
		.mem_outb(mem_outb[226:227]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[228:229]),
		.mem_outb(mem_outb[228:229]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[230:231]),
		.mem_outb(mem_outb[230:231]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[232:233]),
		.mem_outb(mem_outb[232:233]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[234:235]),
		.mem_outb(mem_outb[234:235]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[236:237]),
		.mem_outb(mem_outb[236:237]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[238:239]),
		.mem_outb(mem_outb[238:239]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[240:241]),
		.mem_outb(mem_outb[240:241]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[242:243]),
		.mem_outb(mem_outb[242:243]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[244:245]),
		.mem_outb(mem_outb[244:245]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[246:247]),
		.mem_outb(mem_outb[246:247]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[248:249]),
		.mem_outb(mem_outb[248:249]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[250:251]),
		.mem_outb(mem_outb[250:251]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[252:253]),
		.mem_outb(mem_outb[252:253]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[254:255]),
		.mem_outb(mem_outb[254:255]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[256:257]),
		.mem_outb(mem_outb[256:257]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[258:259]),
		.mem_outb(mem_outb[258:259]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[260:261]),
		.mem_outb(mem_outb[260:261]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[262:263]),
		.mem_outb(mem_outb[262:263]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[264:265]),
		.mem_outb(mem_outb[264:265]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[266:267]),
		.mem_outb(mem_outb[266:267]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[268:269]),
		.mem_outb(mem_outb[268:269]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[270:271]),
		.mem_outb(mem_outb[270:271]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[272:273]),
		.mem_outb(mem_outb[272:273]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[274:275]),
		.mem_outb(mem_outb[274:275]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[276:277]),
		.mem_outb(mem_outb[276:277]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[278:279]),
		.mem_outb(mem_outb[278:279]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[280:281]),
		.mem_outb(mem_outb[280:281]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[282:283]),
		.mem_outb(mem_outb[282:283]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[284:285]),
		.mem_outb(mem_outb[284:285]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[286:287]),
		.mem_outb(mem_outb[286:287]));

	sb_mux_size6_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_0_ccff_tail),
		.mem_out(mem_out[136:138]),
		.mem_outb(mem_outb[136:138]));

	sb_mux_size6_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_1_ccff_tail),
		.mem_out(mem_out[139:141]),
		.mem_outb(mem_outb[139:141]));

	sb_mux_size6_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_2_ccff_tail),
		.mem_out(mem_out[162:164]),
		.mem_outb(mem_outb[162:164]));

	sb_mux_size6_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_3_ccff_tail),
		.mem_out(mem_out[165:167]),
		.mem_outb(mem_outb[165:167]));

	sb_mux_size6_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_4_ccff_tail),
		.mem_out(mem_out[304:306]),
		.mem_outb(mem_outb[304:306]));

	sb_mux_size6_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_5_ccff_tail),
		.mem_out(mem_out[307:309]),
		.mem_outb(mem_outb[307:309]));

	sb_mux_size6_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_6_ccff_tail),
		.mem_out(mem_out[330:332]),
		.mem_outb(mem_outb[330:332]));

	sb_mux_size6_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[333:335]),
		.mem_outb(mem_outb[333:335]));

	sb_mux_size7_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_0_ccff_tail),
		.mem_out(mem_out[150:152]),
		.mem_outb(mem_outb[150:152]));

	sb_mux_size7_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_1_ccff_tail),
		.mem_out(mem_out[153:155]),
		.mem_outb(mem_outb[153:155]));

	sb_mux_size7_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_2_ccff_tail),
		.mem_out(mem_out[156:158]),
		.mem_outb(mem_outb[156:158]));

	sb_mux_size7_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_3_ccff_tail),
		.mem_out(mem_out[159:161]),
		.mem_outb(mem_outb[159:161]));

	sb_mux_size7_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_4_ccff_tail),
		.mem_out(mem_out[318:320]),
		.mem_outb(mem_outb[318:320]));

	sb_mux_size7_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_5_ccff_tail),
		.mem_out(mem_out[321:323]),
		.mem_outb(mem_outb[321:323]));

	sb_mux_size7_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_6_ccff_tail),
		.mem_out(mem_out[324:326]),
		.mem_outb(mem_outb[324:326]));

	sb_mux_size7_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_7_ccff_tail),
		.mem_out(mem_out[327:329]),
		.mem_outb(mem_outb[327:329]));

endmodule
// ----- END Verilog module for sb_10__config_group_mem_size336 -----




// ----- Verilog module for sb_11__config_group_mem_size358 -----
module sb_11__config_group_mem_size358(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:357] mem_out;
//----- OUTPUT PORTS -----
output [0:357] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size15_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size15_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size15_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	sb_mux_size15_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	sb_mux_size15_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_3_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	sb_mux_size15_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size19_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_4_ccff_tail),
		.mem_out(mem_out[39:42]),
		.mem_outb(mem_outb[39:42]));

	sb_mux_size15_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_5_ccff_tail),
		.mem_out(mem_out[43:46]),
		.mem_outb(mem_outb[43:46]));

	sb_mux_size15_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_6_ccff_tail),
		.mem_out(mem_out[47:50]),
		.mem_outb(mem_outb[47:50]));

	sb_mux_size15_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_7_ccff_tail),
		.mem_out(mem_out[179:182]),
		.mem_outb(mem_outb[179:182]));

	sb_mux_size15_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_8_ccff_tail),
		.mem_out(mem_out[183:186]),
		.mem_outb(mem_outb[183:186]));

	sb_mux_size15_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_9_ccff_tail),
		.mem_out(mem_out[187:190]),
		.mem_outb(mem_outb[187:190]));

	sb_mux_size15_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_10_ccff_tail),
		.mem_out(mem_out[191:194]),
		.mem_outb(mem_outb[191:194]));

	sb_mux_size15_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size19_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_11_ccff_tail),
		.mem_out(mem_out[218:221]),
		.mem_outb(mem_outb[218:221]));

	sb_mux_size15_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_12_ccff_tail),
		.mem_out(mem_out[222:225]),
		.mem_outb(mem_outb[222:225]));

	sb_mux_size15_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size15_mem_13_ccff_tail),
		.mem_out(mem_out[226:229]),
		.mem_outb(mem_outb[226:229]));

	sb_mux_size13_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_0_ccff_tail),
		.mem_out(mem_out[16:19]),
		.mem_outb(mem_outb[16:19]));

	sb_mux_size13_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_1_ccff_tail),
		.mem_out(mem_out[51:54]),
		.mem_outb(mem_outb[51:54]));

	sb_mux_size13_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_2_ccff_tail),
		.mem_out(mem_out[55:58]),
		.mem_outb(mem_outb[55:58]));

	sb_mux_size13_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_3_ccff_tail),
		.mem_out(mem_out[195:198]),
		.mem_outb(mem_outb[195:198]));

	sb_mux_size13_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size15_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_4_ccff_tail),
		.mem_out(mem_out[230:233]),
		.mem_outb(mem_outb[230:233]));

	sb_mux_size13_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size13_mem_5_ccff_tail),
		.mem_out(mem_out[234:237]),
		.mem_outb(mem_outb[234:237]));

	sb_mux_size11_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[20:23]),
		.mem_outb(mem_outb[20:23]));

	sb_mux_size11_mem mem_right_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[147:150]),
		.mem_outb(mem_outb[147:150]));

	sb_mux_size11_mem mem_right_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[151:154]),
		.mem_outb(mem_outb[151:154]));

	sb_mux_size11_mem mem_right_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[155:158]),
		.mem_outb(mem_outb[155:158]));

	sb_mux_size11_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_4_ccff_tail),
		.mem_out(mem_out[199:202]),
		.mem_outb(mem_outb[199:202]));

	sb_mux_size11_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_5_ccff_tail),
		.mem_out(mem_out[326:329]),
		.mem_outb(mem_outb[326:329]));

	sb_mux_size11_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_6_ccff_tail),
		.mem_out(mem_out[330:333]),
		.mem_outb(mem_outb[330:333]));

	sb_mux_size11_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_7_ccff_tail),
		.mem_out(mem_out[334:337]),
		.mem_outb(mem_outb[334:337]));

	sb_mux_size21_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size21_mem_0_ccff_tail),
		.mem_out(mem_out[24:28]),
		.mem_outb(mem_outb[24:28]));

	sb_mux_size21_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size21_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size21_mem_1_ccff_tail),
		.mem_out(mem_out[29:33]),
		.mem_outb(mem_outb[29:33]));

	sb_mux_size21_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size21_mem_2_ccff_tail),
		.mem_out(mem_out[203:207]),
		.mem_outb(mem_outb[203:207]));

	sb_mux_size21_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size21_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size21_mem_3_ccff_tail),
		.mem_out(mem_out[208:212]),
		.mem_outb(mem_outb[208:212]));

	sb_mux_size19_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size21_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size19_mem_0_ccff_tail),
		.mem_out(mem_out[34:38]),
		.mem_outb(mem_outb[34:38]));

	sb_mux_size19_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size21_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size19_mem_1_ccff_tail),
		.mem_out(mem_out[213:217]),
		.mem_outb(mem_outb[213:217]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[59:60]),
		.mem_outb(mem_outb[59:60]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[61:62]),
		.mem_outb(mem_outb[61:62]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[63:64]),
		.mem_outb(mem_outb[63:64]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[65:66]),
		.mem_outb(mem_outb[65:66]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[67:68]),
		.mem_outb(mem_outb[67:68]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[69:70]),
		.mem_outb(mem_outb[69:70]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[71:72]),
		.mem_outb(mem_outb[71:72]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[73:74]),
		.mem_outb(mem_outb[73:74]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[75:76]),
		.mem_outb(mem_outb[75:76]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[77:78]),
		.mem_outb(mem_outb[77:78]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[79:80]),
		.mem_outb(mem_outb[79:80]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[81:82]),
		.mem_outb(mem_outb[81:82]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[83:84]),
		.mem_outb(mem_outb[83:84]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[85:86]),
		.mem_outb(mem_outb[85:86]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[87:88]),
		.mem_outb(mem_outb[87:88]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[89:90]),
		.mem_outb(mem_outb[89:90]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[91:92]),
		.mem_outb(mem_outb[91:92]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[93:94]),
		.mem_outb(mem_outb[93:94]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[95:96]),
		.mem_outb(mem_outb[95:96]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[97:98]),
		.mem_outb(mem_outb[97:98]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[99:100]),
		.mem_outb(mem_outb[99:100]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[101:102]),
		.mem_outb(mem_outb[101:102]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[103:104]),
		.mem_outb(mem_outb[103:104]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[105:106]),
		.mem_outb(mem_outb[105:106]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[107:108]),
		.mem_outb(mem_outb[107:108]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[109:110]),
		.mem_outb(mem_outb[109:110]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[111:112]),
		.mem_outb(mem_outb[111:112]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[113:114]),
		.mem_outb(mem_outb[113:114]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[115:116]),
		.mem_outb(mem_outb[115:116]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[117:118]),
		.mem_outb(mem_outb[117:118]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[119:120]),
		.mem_outb(mem_outb[119:120]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[121:122]),
		.mem_outb(mem_outb[121:122]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size13_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[238:239]),
		.mem_outb(mem_outb[238:239]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[240:241]),
		.mem_outb(mem_outb[240:241]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[242:243]),
		.mem_outb(mem_outb[242:243]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[244:245]),
		.mem_outb(mem_outb[244:245]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[246:247]),
		.mem_outb(mem_outb[246:247]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[248:249]),
		.mem_outb(mem_outb[248:249]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[250:251]),
		.mem_outb(mem_outb[250:251]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[252:253]),
		.mem_outb(mem_outb[252:253]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[254:255]),
		.mem_outb(mem_outb[254:255]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[256:257]),
		.mem_outb(mem_outb[256:257]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[258:259]),
		.mem_outb(mem_outb[258:259]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[260:261]),
		.mem_outb(mem_outb[260:261]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[262:263]),
		.mem_outb(mem_outb[262:263]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[264:265]),
		.mem_outb(mem_outb[264:265]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[266:267]),
		.mem_outb(mem_outb[266:267]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[268:269]),
		.mem_outb(mem_outb[268:269]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[270:271]),
		.mem_outb(mem_outb[270:271]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[272:273]),
		.mem_outb(mem_outb[272:273]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[274:275]),
		.mem_outb(mem_outb[274:275]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[276:277]),
		.mem_outb(mem_outb[276:277]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[278:279]),
		.mem_outb(mem_outb[278:279]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[280:281]),
		.mem_outb(mem_outb[280:281]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[282:283]),
		.mem_outb(mem_outb[282:283]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[284:285]),
		.mem_outb(mem_outb[284:285]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[286:287]),
		.mem_outb(mem_outb[286:287]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[288:289]),
		.mem_outb(mem_outb[288:289]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[290:291]),
		.mem_outb(mem_outb[290:291]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[292:293]),
		.mem_outb(mem_outb[292:293]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[294:295]),
		.mem_outb(mem_outb[294:295]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[296:297]),
		.mem_outb(mem_outb[296:297]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[298:299]),
		.mem_outb(mem_outb[298:299]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[300:301]),
		.mem_outb(mem_outb[300:301]));

	sb_mux_size10_mem mem_right_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[123:126]),
		.mem_outb(mem_outb[123:126]));

	sb_mux_size10_mem mem_right_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[127:130]),
		.mem_outb(mem_outb[127:130]));

	sb_mux_size10_mem mem_right_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_2_ccff_tail),
		.mem_out(mem_out[131:134]),
		.mem_outb(mem_outb[131:134]));

	sb_mux_size10_mem mem_right_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_3_ccff_tail),
		.mem_out(mem_out[135:138]),
		.mem_outb(mem_outb[135:138]));

	sb_mux_size10_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_4_ccff_tail),
		.mem_out(mem_out[302:305]),
		.mem_outb(mem_outb[302:305]));

	sb_mux_size10_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_5_ccff_tail),
		.mem_out(mem_out[306:309]),
		.mem_outb(mem_outb[306:309]));

	sb_mux_size10_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_6_ccff_tail),
		.mem_out(mem_out[310:313]),
		.mem_outb(mem_outb[310:313]));

	sb_mux_size10_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_7_ccff_tail),
		.mem_out(mem_out[314:317]),
		.mem_outb(mem_outb[314:317]));

	sb_mux_size8_mem mem_right_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[139:142]),
		.mem_outb(mem_outb[139:142]));

	sb_mux_size8_mem mem_right_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[143:146]),
		.mem_outb(mem_outb[143:146]));

	sb_mux_size8_mem mem_right_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[171:174]),
		.mem_outb(mem_outb[171:174]));

	sb_mux_size8_mem mem_right_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[175:178]),
		.mem_outb(mem_outb[175:178]));

	sb_mux_size8_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[318:321]),
		.mem_outb(mem_outb[318:321]));

	sb_mux_size8_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[322:325]),
		.mem_outb(mem_outb[322:325]));

	sb_mux_size8_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[350:353]),
		.mem_outb(mem_outb[350:353]));

	sb_mux_size8_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[354:357]),
		.mem_outb(mem_outb[354:357]));

	sb_mux_size9_mem mem_right_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[159:162]),
		.mem_outb(mem_outb[159:162]));

	sb_mux_size9_mem mem_right_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_1_ccff_tail),
		.mem_out(mem_out[163:166]),
		.mem_outb(mem_outb[163:166]));

	sb_mux_size9_mem mem_right_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_2_ccff_tail),
		.mem_out(mem_out[167:170]),
		.mem_outb(mem_outb[167:170]));

	sb_mux_size9_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_3_ccff_tail),
		.mem_out(mem_out[338:341]),
		.mem_outb(mem_outb[338:341]));

	sb_mux_size9_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_4_ccff_tail),
		.mem_out(mem_out[342:345]),
		.mem_outb(mem_outb[342:345]));

	sb_mux_size9_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_5_ccff_tail),
		.mem_out(mem_out[346:349]),
		.mem_outb(mem_outb[346:349]));

endmodule
// ----- END Verilog module for sb_11__config_group_mem_size358 -----




// ----- Verilog module for sb_12__config_group_mem_size315 -----
module sb_12__config_group_mem_size315(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:314] mem_out;
//----- OUTPUT PORTS -----
output [0:314] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size8_mem mem_top_track_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(sb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	sb_mux_size8_mem mem_top_track_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[31:34]),
		.mem_outb(mem_outb[31:34]));

	sb_mux_size8_mem mem_top_track_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[35:38]),
		.mem_outb(mem_outb[35:38]));

	sb_mux_size8_mem mem_top_track_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size9_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[43:46]),
		.mem_outb(mem_outb[43:46]));

	sb_mux_size8_mem mem_top_track_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[47:50]),
		.mem_outb(mem_outb[47:50]));

	sb_mux_size8_mem mem_bottom_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_31_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[115:118]),
		.mem_outb(mem_outb[115:118]));

	sb_mux_size8_mem mem_bottom_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[119:122]),
		.mem_outb(mem_outb[119:122]));

	sb_mux_size8_mem mem_bottom_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[123:126]),
		.mem_outb(mem_outb[123:126]));

	sb_mux_size8_mem mem_bottom_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size10_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[148:151]),
		.mem_outb(mem_outb[148:151]));

	sb_mux_size8_mem mem_bottom_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[152:155]),
		.mem_outb(mem_outb[152:155]));

	sb_mux_size8_mem mem_bottom_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_10_ccff_tail),
		.mem_out(mem_out[156:159]),
		.mem_outb(mem_outb[156:159]));

	sb_mux_size8_mem mem_bottom_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_11_ccff_tail),
		.mem_out(mem_out[163:166]),
		.mem_outb(mem_outb[163:166]));

	sb_mux_size8_mem mem_left_track_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_63_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_12_ccff_tail),
		.mem_out(mem_out[231:234]),
		.mem_outb(mem_outb[231:234]));

	sb_mux_size8_mem mem_left_track_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_13_ccff_tail),
		.mem_out(mem_out[235:238]),
		.mem_outb(mem_outb[235:238]));

	sb_mux_size8_mem mem_left_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_14_ccff_tail),
		.mem_out(mem_out[251:254]),
		.mem_outb(mem_outb[251:254]));

	sb_mux_size8_mem mem_left_track_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size8_mem_15_ccff_tail),
		.mem_out(mem_out[255:258]),
		.mem_outb(mem_outb[255:258]));

	sb_mux_size7_mem mem_top_track_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_0_ccff_tail),
		.mem_out(mem_out[4:6]),
		.mem_outb(mem_outb[4:6]));

	sb_mux_size7_mem mem_top_track_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_1_ccff_tail),
		.mem_out(mem_out[7:9]),
		.mem_outb(mem_outb[7:9]));

	sb_mux_size7_mem mem_top_track_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_2_ccff_tail),
		.mem_out(mem_out[10:12]),
		.mem_outb(mem_outb[10:12]));

	sb_mux_size7_mem mem_top_track_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_3_ccff_tail),
		.mem_out(mem_out[13:15]),
		.mem_outb(mem_outb[13:15]));

	sb_mux_size7_mem mem_bottom_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_4_ccff_tail),
		.mem_out(mem_out[127:129]),
		.mem_outb(mem_outb[127:129]));

	sb_mux_size7_mem mem_bottom_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_5_ccff_tail),
		.mem_out(mem_out[130:132]),
		.mem_outb(mem_outb[130:132]));

	sb_mux_size7_mem mem_bottom_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_6_ccff_tail),
		.mem_out(mem_out[160:162]),
		.mem_outb(mem_outb[160:162]));

	sb_mux_size7_mem mem_left_track_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_7_ccff_tail),
		.mem_out(mem_out[239:241]),
		.mem_outb(mem_outb[239:241]));

	sb_mux_size7_mem mem_left_track_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_8_ccff_tail),
		.mem_out(mem_out[242:244]),
		.mem_outb(mem_outb[242:244]));

	sb_mux_size7_mem mem_left_track_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_9_ccff_tail),
		.mem_out(mem_out[245:247]),
		.mem_outb(mem_outb[245:247]));

	sb_mux_size7_mem mem_left_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_10_ccff_tail),
		.mem_out(mem_out[248:250]),
		.mem_outb(mem_outb[248:250]));

	sb_mux_size7_mem mem_left_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_15_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_11_ccff_tail),
		.mem_out(mem_out[259:261]),
		.mem_outb(mem_outb[259:261]));

	sb_mux_size7_mem mem_left_track_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_11_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_12_ccff_tail),
		.mem_out(mem_out[262:264]),
		.mem_outb(mem_outb[262:264]));

	sb_mux_size7_mem mem_left_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_12_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_13_ccff_tail),
		.mem_out(mem_out[265:267]),
		.mem_outb(mem_outb[265:267]));

	sb_mux_size7_mem mem_left_track_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_13_ccff_tail),
		.ccff_tail(sb_mux_size7_mem_14_ccff_tail),
		.mem_out(mem_out[268:270]),
		.mem_outb(mem_outb[268:270]));

	sb_mux_size6_mem mem_top_track_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_0_ccff_tail),
		.mem_out(mem_out[16:18]),
		.mem_outb(mem_outb[16:18]));

	sb_mux_size6_mem mem_bottom_track_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size6_mem_1_ccff_tail),
		.mem_out(mem_out[133:135]),
		.mem_outb(mem_outb[133:135]));

	sb_mux_size11_mem mem_top_track_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_0_ccff_tail),
		.mem_out(mem_out[19:22]),
		.mem_outb(mem_outb[19:22]));

	sb_mux_size11_mem mem_top_track_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_1_ccff_tail),
		.mem_out(mem_out[23:26]),
		.mem_outb(mem_outb[23:26]));

	sb_mux_size11_mem mem_bottom_track_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size6_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_2_ccff_tail),
		.mem_out(mem_out[136:139]),
		.mem_outb(mem_outb[136:139]));

	sb_mux_size11_mem mem_bottom_track_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size11_mem_3_ccff_tail),
		.mem_out(mem_out[140:143]),
		.mem_outb(mem_outb[140:143]));

	sb_mux_size10_mem mem_top_track_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_0_ccff_tail),
		.mem_out(mem_out[27:30]),
		.mem_outb(mem_outb[27:30]));

	sb_mux_size10_mem mem_bottom_track_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size11_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size10_mem_1_ccff_tail),
		.mem_out(mem_out[144:147]),
		.mem_outb(mem_outb[144:147]));

	sb_mux_size9_mem mem_top_track_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size9_mem_0_ccff_tail),
		.mem_out(mem_out[39:42]),
		.mem_outb(mem_outb[39:42]));

	clk_mux_size3_mem mem_top_track_64 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_0_ccff_tail),
		.mem_out(mem_out[51:52]),
		.mem_outb(mem_outb[51:52]));

	clk_mux_size3_mem mem_top_track_66 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_0_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_1_ccff_tail),
		.mem_out(mem_out[53:54]),
		.mem_outb(mem_outb[53:54]));

	clk_mux_size3_mem mem_top_track_68 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_1_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_2_ccff_tail),
		.mem_out(mem_out[55:56]),
		.mem_outb(mem_outb[55:56]));

	clk_mux_size3_mem mem_top_track_70 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_2_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_3_ccff_tail),
		.mem_out(mem_out[57:58]),
		.mem_outb(mem_outb[57:58]));

	clk_mux_size3_mem mem_top_track_72 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_3_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_4_ccff_tail),
		.mem_out(mem_out[59:60]),
		.mem_outb(mem_outb[59:60]));

	clk_mux_size3_mem mem_top_track_74 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_4_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_5_ccff_tail),
		.mem_out(mem_out[61:62]),
		.mem_outb(mem_outb[61:62]));

	clk_mux_size3_mem mem_top_track_76 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_5_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_6_ccff_tail),
		.mem_out(mem_out[63:64]),
		.mem_outb(mem_outb[63:64]));

	clk_mux_size3_mem mem_top_track_78 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_6_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_7_ccff_tail),
		.mem_out(mem_out[65:66]),
		.mem_outb(mem_outb[65:66]));

	clk_mux_size3_mem mem_top_track_80 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_7_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_8_ccff_tail),
		.mem_out(mem_out[67:68]),
		.mem_outb(mem_outb[67:68]));

	clk_mux_size3_mem mem_top_track_82 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_8_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_9_ccff_tail),
		.mem_out(mem_out[69:70]),
		.mem_outb(mem_outb[69:70]));

	clk_mux_size3_mem mem_top_track_84 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_9_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_10_ccff_tail),
		.mem_out(mem_out[71:72]),
		.mem_outb(mem_outb[71:72]));

	clk_mux_size3_mem mem_top_track_86 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_10_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_11_ccff_tail),
		.mem_out(mem_out[73:74]),
		.mem_outb(mem_outb[73:74]));

	clk_mux_size3_mem mem_top_track_88 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_12_ccff_tail),
		.mem_out(mem_out[75:76]),
		.mem_outb(mem_outb[75:76]));

	clk_mux_size3_mem mem_top_track_90 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_12_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_13_ccff_tail),
		.mem_out(mem_out[77:78]),
		.mem_outb(mem_outb[77:78]));

	clk_mux_size3_mem mem_top_track_92 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_13_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_14_ccff_tail),
		.mem_out(mem_out[79:80]),
		.mem_outb(mem_outb[79:80]));

	clk_mux_size3_mem mem_top_track_94 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_14_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_15_ccff_tail),
		.mem_out(mem_out[81:82]),
		.mem_outb(mem_outb[81:82]));

	clk_mux_size3_mem mem_top_track_96 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_15_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_16_ccff_tail),
		.mem_out(mem_out[83:84]),
		.mem_outb(mem_outb[83:84]));

	clk_mux_size3_mem mem_top_track_98 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_16_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_17_ccff_tail),
		.mem_out(mem_out[85:86]),
		.mem_outb(mem_outb[85:86]));

	clk_mux_size3_mem mem_top_track_100 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_17_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_18_ccff_tail),
		.mem_out(mem_out[87:88]),
		.mem_outb(mem_outb[87:88]));

	clk_mux_size3_mem mem_top_track_102 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_18_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_19_ccff_tail),
		.mem_out(mem_out[89:90]),
		.mem_outb(mem_outb[89:90]));

	clk_mux_size3_mem mem_top_track_104 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_19_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_20_ccff_tail),
		.mem_out(mem_out[91:92]),
		.mem_outb(mem_outb[91:92]));

	clk_mux_size3_mem mem_top_track_106 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_20_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_21_ccff_tail),
		.mem_out(mem_out[93:94]),
		.mem_outb(mem_outb[93:94]));

	clk_mux_size3_mem mem_top_track_108 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_21_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_22_ccff_tail),
		.mem_out(mem_out[95:96]),
		.mem_outb(mem_outb[95:96]));

	clk_mux_size3_mem mem_top_track_110 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_22_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_23_ccff_tail),
		.mem_out(mem_out[97:98]),
		.mem_outb(mem_outb[97:98]));

	clk_mux_size3_mem mem_top_track_112 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_23_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_24_ccff_tail),
		.mem_out(mem_out[99:100]),
		.mem_outb(mem_outb[99:100]));

	clk_mux_size3_mem mem_top_track_114 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_24_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_25_ccff_tail),
		.mem_out(mem_out[101:102]),
		.mem_outb(mem_outb[101:102]));

	clk_mux_size3_mem mem_top_track_116 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_25_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_26_ccff_tail),
		.mem_out(mem_out[103:104]),
		.mem_outb(mem_outb[103:104]));

	clk_mux_size3_mem mem_top_track_118 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_26_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_27_ccff_tail),
		.mem_out(mem_out[105:106]),
		.mem_outb(mem_outb[105:106]));

	clk_mux_size3_mem mem_top_track_120 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_27_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_28_ccff_tail),
		.mem_out(mem_out[107:108]),
		.mem_outb(mem_outb[107:108]));

	clk_mux_size3_mem mem_top_track_122 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_28_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_29_ccff_tail),
		.mem_out(mem_out[109:110]),
		.mem_outb(mem_outb[109:110]));

	clk_mux_size3_mem mem_top_track_124 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_29_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_30_ccff_tail),
		.mem_out(mem_out[111:112]),
		.mem_outb(mem_outb[111:112]));

	clk_mux_size3_mem mem_top_track_126 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_30_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_31_ccff_tail),
		.mem_out(mem_out[113:114]),
		.mem_outb(mem_outb[113:114]));

	clk_mux_size3_mem mem_bottom_track_65 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size8_mem_11_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_32_ccff_tail),
		.mem_out(mem_out[167:168]),
		.mem_outb(mem_outb[167:168]));

	clk_mux_size3_mem mem_bottom_track_67 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_32_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_33_ccff_tail),
		.mem_out(mem_out[169:170]),
		.mem_outb(mem_outb[169:170]));

	clk_mux_size3_mem mem_bottom_track_69 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_33_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_34_ccff_tail),
		.mem_out(mem_out[171:172]),
		.mem_outb(mem_outb[171:172]));

	clk_mux_size3_mem mem_bottom_track_71 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_34_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_35_ccff_tail),
		.mem_out(mem_out[173:174]),
		.mem_outb(mem_outb[173:174]));

	clk_mux_size3_mem mem_bottom_track_73 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_35_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_36_ccff_tail),
		.mem_out(mem_out[175:176]),
		.mem_outb(mem_outb[175:176]));

	clk_mux_size3_mem mem_bottom_track_75 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_36_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_37_ccff_tail),
		.mem_out(mem_out[177:178]),
		.mem_outb(mem_outb[177:178]));

	clk_mux_size3_mem mem_bottom_track_77 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_37_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_38_ccff_tail),
		.mem_out(mem_out[179:180]),
		.mem_outb(mem_outb[179:180]));

	clk_mux_size3_mem mem_bottom_track_79 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_38_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_39_ccff_tail),
		.mem_out(mem_out[181:182]),
		.mem_outb(mem_outb[181:182]));

	clk_mux_size3_mem mem_bottom_track_81 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_39_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_40_ccff_tail),
		.mem_out(mem_out[183:184]),
		.mem_outb(mem_outb[183:184]));

	clk_mux_size3_mem mem_bottom_track_83 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_40_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_41_ccff_tail),
		.mem_out(mem_out[185:186]),
		.mem_outb(mem_outb[185:186]));

	clk_mux_size3_mem mem_bottom_track_85 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_41_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_42_ccff_tail),
		.mem_out(mem_out[187:188]),
		.mem_outb(mem_outb[187:188]));

	clk_mux_size3_mem mem_bottom_track_87 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_42_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_43_ccff_tail),
		.mem_out(mem_out[189:190]),
		.mem_outb(mem_outb[189:190]));

	clk_mux_size3_mem mem_bottom_track_89 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_43_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_44_ccff_tail),
		.mem_out(mem_out[191:192]),
		.mem_outb(mem_outb[191:192]));

	clk_mux_size3_mem mem_bottom_track_91 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_44_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_45_ccff_tail),
		.mem_out(mem_out[193:194]),
		.mem_outb(mem_outb[193:194]));

	clk_mux_size3_mem mem_bottom_track_93 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_45_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_46_ccff_tail),
		.mem_out(mem_out[195:196]),
		.mem_outb(mem_outb[195:196]));

	clk_mux_size3_mem mem_bottom_track_95 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_46_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_47_ccff_tail),
		.mem_out(mem_out[197:198]),
		.mem_outb(mem_outb[197:198]));

	clk_mux_size3_mem mem_bottom_track_97 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_47_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_48_ccff_tail),
		.mem_out(mem_out[199:200]),
		.mem_outb(mem_outb[199:200]));

	clk_mux_size3_mem mem_bottom_track_99 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_48_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_49_ccff_tail),
		.mem_out(mem_out[201:202]),
		.mem_outb(mem_outb[201:202]));

	clk_mux_size3_mem mem_bottom_track_101 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_49_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_50_ccff_tail),
		.mem_out(mem_out[203:204]),
		.mem_outb(mem_outb[203:204]));

	clk_mux_size3_mem mem_bottom_track_103 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_50_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_51_ccff_tail),
		.mem_out(mem_out[205:206]),
		.mem_outb(mem_outb[205:206]));

	clk_mux_size3_mem mem_bottom_track_105 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_51_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_52_ccff_tail),
		.mem_out(mem_out[207:208]),
		.mem_outb(mem_outb[207:208]));

	clk_mux_size3_mem mem_bottom_track_107 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_52_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_53_ccff_tail),
		.mem_out(mem_out[209:210]),
		.mem_outb(mem_outb[209:210]));

	clk_mux_size3_mem mem_bottom_track_109 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_53_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_54_ccff_tail),
		.mem_out(mem_out[211:212]),
		.mem_outb(mem_outb[211:212]));

	clk_mux_size3_mem mem_bottom_track_111 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_54_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_55_ccff_tail),
		.mem_out(mem_out[213:214]),
		.mem_outb(mem_outb[213:214]));

	clk_mux_size3_mem mem_bottom_track_113 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_55_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_56_ccff_tail),
		.mem_out(mem_out[215:216]),
		.mem_outb(mem_outb[215:216]));

	clk_mux_size3_mem mem_bottom_track_115 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_56_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_57_ccff_tail),
		.mem_out(mem_out[217:218]),
		.mem_outb(mem_outb[217:218]));

	clk_mux_size3_mem mem_bottom_track_117 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_57_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_58_ccff_tail),
		.mem_out(mem_out[219:220]),
		.mem_outb(mem_outb[219:220]));

	clk_mux_size3_mem mem_bottom_track_119 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_58_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_59_ccff_tail),
		.mem_out(mem_out[221:222]),
		.mem_outb(mem_outb[221:222]));

	clk_mux_size3_mem mem_bottom_track_121 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_59_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_60_ccff_tail),
		.mem_out(mem_out[223:224]),
		.mem_outb(mem_outb[223:224]));

	clk_mux_size3_mem mem_bottom_track_123 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_60_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_61_ccff_tail),
		.mem_out(mem_out[225:226]),
		.mem_outb(mem_outb[225:226]));

	clk_mux_size3_mem mem_bottom_track_125 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_61_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_62_ccff_tail),
		.mem_out(mem_out[227:228]),
		.mem_outb(mem_outb[227:228]));

	clk_mux_size3_mem mem_bottom_track_127 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(clk_mux_size3_mem_62_ccff_tail),
		.ccff_tail(clk_mux_size3_mem_63_ccff_tail),
		.mem_out(mem_out[229:230]),
		.mem_outb(mem_outb[229:230]));

	sb_mux_size5_mem mem_left_track_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size7_mem_14_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_0_ccff_tail),
		.mem_out(mem_out[271:273]),
		.mem_outb(mem_outb[271:273]));

	sb_mux_size5_mem mem_left_track_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_1_ccff_tail),
		.mem_out(mem_out[274:276]),
		.mem_outb(mem_outb[274:276]));

	sb_mux_size5_mem mem_left_track_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size5_mem_2_ccff_tail),
		.mem_out(mem_out[277:279]),
		.mem_outb(mem_outb[277:279]));

	sb_mux_size4_mem mem_left_track_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size5_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_0_ccff_tail),
		.mem_out(mem_out[280:282]),
		.mem_outb(mem_outb[280:282]));

	sb_mux_size4_mem mem_left_track_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_1_ccff_tail),
		.mem_out(mem_out[283:285]),
		.mem_outb(mem_outb[283:285]));

	sb_mux_size4_mem mem_left_track_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size4_mem_2_ccff_tail),
		.mem_out(mem_out[286:288]),
		.mem_outb(mem_outb[286:288]));

	sb_mux_size2_mem mem_left_track_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size4_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_0_ccff_tail),
		.mem_out(mem_out[289:290]),
		.mem_outb(mem_outb[289:290]));

	sb_mux_size2_mem mem_left_track_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_0_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_1_ccff_tail),
		.mem_out(mem_out[291:292]),
		.mem_outb(mem_outb[291:292]));

	sb_mux_size2_mem mem_left_track_43 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_1_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_2_ccff_tail),
		.mem_out(mem_out[293:294]),
		.mem_outb(mem_outb[293:294]));

	sb_mux_size2_mem mem_left_track_45 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_2_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_3_ccff_tail),
		.mem_out(mem_out[295:296]),
		.mem_outb(mem_outb[295:296]));

	sb_mux_size2_mem mem_left_track_47 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_3_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_4_ccff_tail),
		.mem_out(mem_out[297:298]),
		.mem_outb(mem_outb[297:298]));

	sb_mux_size2_mem mem_left_track_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_4_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_5_ccff_tail),
		.mem_out(mem_out[299:300]),
		.mem_outb(mem_outb[299:300]));

	sb_mux_size2_mem mem_left_track_51 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_5_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_6_ccff_tail),
		.mem_out(mem_out[301:302]),
		.mem_outb(mem_outb[301:302]));

	sb_mux_size2_mem mem_left_track_53 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_6_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_7_ccff_tail),
		.mem_out(mem_out[303:304]),
		.mem_outb(mem_outb[303:304]));

	sb_mux_size2_mem mem_left_track_55 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_7_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_8_ccff_tail),
		.mem_out(mem_out[305:306]),
		.mem_outb(mem_outb[305:306]));

	sb_mux_size2_mem mem_left_track_57 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_8_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_9_ccff_tail),
		.mem_out(mem_out[307:308]),
		.mem_outb(mem_outb[307:308]));

	sb_mux_size2_mem mem_left_track_59 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_9_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_10_ccff_tail),
		.mem_out(mem_out[309:310]),
		.mem_outb(mem_outb[309:310]));

	sb_mux_size2_mem mem_left_track_61 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_10_ccff_tail),
		.ccff_tail(sb_mux_size2_mem_11_ccff_tail),
		.mem_out(mem_out[311:312]),
		.mem_outb(mem_outb[311:312]));

	sb_mux_size2_mem mem_left_track_63 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(sb_mux_size2_mem_11_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[313:314]),
		.mem_outb(mem_outb[313:314]));

endmodule
// ----- END Verilog module for sb_12__config_group_mem_size315 -----




// ----- Verilog module for cbx_2__config_group_mem_size32 -----
module cbx_2__config_group_mem_size32(config_enable,
                                      prog_reset,
                                      prog_clk,
                                      ccff_head,
                                      mem_out,
                                      mem_outb,
                                      ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:31] mem_out;
//----- OUTPUT PORTS -----
output [0:31] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size8_mem mem_top_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	cb_mux_size8_mem mem_top_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	cb_mux_size8_mem mem_top_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	cb_mux_size8_mem mem_top_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	cb_mux_size8_mem mem_top_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[16:19]),
		.mem_outb(mem_outb[16:19]));

	cb_mux_size8_mem mem_top_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[20:23]),
		.mem_outb(mem_outb[20:23]));

	cb_mux_size8_mem mem_top_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[24:27]),
		.mem_outb(mem_outb[24:27]));

	cb_mux_size8_mem mem_top_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[28:31]),
		.mem_outb(mem_outb[28:31]));

endmodule
// ----- END Verilog module for cbx_2__config_group_mem_size32 -----




// ----- Verilog module for cbx_3__config_group_mem_size174 -----
module cbx_3__config_group_mem_size174(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:173] mem_out;
//----- OUTPUT PORTS -----
output [0:173] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size26_mem mem_top_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size26_mem_0_ccff_tail),
		.mem_out(mem_out[0:4]),
		.mem_outb(mem_outb[0:4]));

	cb_mux_size26_mem mem_top_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_1_ccff_tail),
		.mem_out(mem_out[5:9]),
		.mem_outb(mem_outb[5:9]));

	cb_mux_size26_mem mem_top_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_2_ccff_tail),
		.mem_out(mem_out[10:14]),
		.mem_outb(mem_outb[10:14]));

	cb_mux_size26_mem mem_top_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_3_ccff_tail),
		.mem_out(mem_out[15:19]),
		.mem_outb(mem_outb[15:19]));

	cb_mux_size26_mem mem_top_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_4_ccff_tail),
		.mem_out(mem_out[20:24]),
		.mem_outb(mem_outb[20:24]));

	cb_mux_size26_mem mem_top_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_5_ccff_tail),
		.mem_out(mem_out[25:29]),
		.mem_outb(mem_outb[25:29]));

	cb_mux_size26_mem mem_top_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_6_ccff_tail),
		.mem_out(mem_out[30:34]),
		.mem_outb(mem_outb[30:34]));

	cb_mux_size26_mem mem_top_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_7_ccff_tail),
		.mem_out(mem_out[35:39]),
		.mem_outb(mem_outb[35:39]));

	cb_mux_size26_mem mem_top_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_8_ccff_tail),
		.mem_out(mem_out[40:44]),
		.mem_outb(mem_outb[40:44]));

	cb_mux_size26_mem mem_top_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_9_ccff_tail),
		.mem_out(mem_out[45:49]),
		.mem_outb(mem_outb[45:49]));

	cb_mux_size26_mem mem_top_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_10_ccff_tail),
		.mem_out(mem_out[50:54]),
		.mem_outb(mem_outb[50:54]));

	cb_mux_size26_mem mem_top_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_11_ccff_tail),
		.mem_out(mem_out[55:59]),
		.mem_outb(mem_outb[55:59]));

	cb_mux_size26_mem mem_top_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_12_ccff_tail),
		.mem_out(mem_out[60:64]),
		.mem_outb(mem_outb[60:64]));

	cb_mux_size26_mem mem_top_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_13_ccff_tail),
		.mem_out(mem_out[65:69]),
		.mem_outb(mem_outb[65:69]));

	cb_mux_size26_mem mem_top_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_14_ccff_tail),
		.mem_out(mem_out[70:74]),
		.mem_outb(mem_outb[70:74]));

	cb_mux_size26_mem mem_top_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_15_ccff_tail),
		.mem_out(mem_out[75:79]),
		.mem_outb(mem_outb[75:79]));

	cb_mux_size26_mem mem_top_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_16_ccff_tail),
		.mem_out(mem_out[80:84]),
		.mem_outb(mem_outb[80:84]));

	cb_mux_size26_mem mem_top_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_17_ccff_tail),
		.mem_out(mem_out[85:89]),
		.mem_outb(mem_outb[85:89]));

	cb_mux_size26_mem mem_top_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_18_ccff_tail),
		.mem_out(mem_out[90:94]),
		.mem_outb(mem_outb[90:94]));

	cb_mux_size26_mem mem_top_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_19_ccff_tail),
		.mem_out(mem_out[95:99]),
		.mem_outb(mem_outb[95:99]));

	cb_mux_size26_mem mem_top_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_20_ccff_tail),
		.mem_out(mem_out[100:104]),
		.mem_outb(mem_outb[100:104]));

	cb_mux_size26_mem mem_top_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_21_ccff_tail),
		.mem_out(mem_out[105:109]),
		.mem_outb(mem_outb[105:109]));

	cb_mux_size26_mem mem_top_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_22_ccff_tail),
		.mem_out(mem_out[110:114]),
		.mem_outb(mem_outb[110:114]));

	cb_mux_size26_mem mem_top_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_23_ccff_tail),
		.mem_out(mem_out[115:119]),
		.mem_outb(mem_outb[115:119]));

	cb_mux_size26_mem mem_top_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_24_ccff_tail),
		.mem_out(mem_out[120:124]),
		.mem_outb(mem_outb[120:124]));

	cb_mux_size26_mem mem_top_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_25_ccff_tail),
		.mem_out(mem_out[125:129]),
		.mem_outb(mem_outb[125:129]));

	cb_mux_size26_mem mem_top_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_26_ccff_tail),
		.mem_out(mem_out[130:134]),
		.mem_outb(mem_outb[130:134]));

	cb_mux_size26_mem mem_top_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_27_ccff_tail),
		.mem_out(mem_out[135:139]),
		.mem_outb(mem_outb[135:139]));

	cb_mux_size26_mem mem_top_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_28_ccff_tail),
		.mem_out(mem_out[140:144]),
		.mem_outb(mem_outb[140:144]));

	cb_mux_size26_mem mem_top_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_29_ccff_tail),
		.mem_out(mem_out[145:149]),
		.mem_outb(mem_outb[145:149]));

	cb_mux_size8_mem mem_top_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[150:153]),
		.mem_outb(mem_outb[150:153]));

	cb_mux_size8_mem mem_top_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[154:157]),
		.mem_outb(mem_outb[154:157]));

	cb_mux_size8_mem mem_top_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[158:161]),
		.mem_outb(mem_outb[158:161]));

	cb_mux_size8_mem mem_top_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[162:165]),
		.mem_outb(mem_outb[162:165]));

	cb_mux_size8_mem mem_top_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[166:169]),
		.mem_outb(mem_outb[166:169]));

	cb_mux_size8_mem mem_top_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[170:173]),
		.mem_outb(mem_outb[170:173]));

endmodule
// ----- END Verilog module for cbx_3__config_group_mem_size174 -----




// ----- Verilog module for cbx_4__config_group_mem_size206 -----
module cbx_4__config_group_mem_size206(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:205] mem_out;
//----- OUTPUT PORTS -----
output [0:205] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size8_mem mem_bottom_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	cb_mux_size8_mem mem_bottom_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	cb_mux_size8_mem mem_bottom_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	cb_mux_size8_mem mem_bottom_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	cb_mux_size8_mem mem_bottom_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[16:19]),
		.mem_outb(mem_outb[16:19]));

	cb_mux_size8_mem mem_bottom_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[20:23]),
		.mem_outb(mem_outb[20:23]));

	cb_mux_size8_mem mem_bottom_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[24:27]),
		.mem_outb(mem_outb[24:27]));

	cb_mux_size8_mem mem_bottom_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[28:31]),
		.mem_outb(mem_outb[28:31]));

	cb_mux_size8_mem mem_top_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[182:185]),
		.mem_outb(mem_outb[182:185]));

	cb_mux_size8_mem mem_top_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[186:189]),
		.mem_outb(mem_outb[186:189]));

	cb_mux_size8_mem mem_top_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_10_ccff_tail),
		.mem_out(mem_out[190:193]),
		.mem_outb(mem_outb[190:193]));

	cb_mux_size8_mem mem_top_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_11_ccff_tail),
		.mem_out(mem_out[194:197]),
		.mem_outb(mem_outb[194:197]));

	cb_mux_size8_mem mem_top_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_12_ccff_tail),
		.mem_out(mem_out[198:201]),
		.mem_outb(mem_outb[198:201]));

	cb_mux_size8_mem mem_top_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_12_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[202:205]),
		.mem_outb(mem_outb[202:205]));

	cb_mux_size26_mem mem_top_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_0_ccff_tail),
		.mem_out(mem_out[32:36]),
		.mem_outb(mem_outb[32:36]));

	cb_mux_size26_mem mem_top_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_1_ccff_tail),
		.mem_out(mem_out[37:41]),
		.mem_outb(mem_outb[37:41]));

	cb_mux_size26_mem mem_top_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_2_ccff_tail),
		.mem_out(mem_out[42:46]),
		.mem_outb(mem_outb[42:46]));

	cb_mux_size26_mem mem_top_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_3_ccff_tail),
		.mem_out(mem_out[47:51]),
		.mem_outb(mem_outb[47:51]));

	cb_mux_size26_mem mem_top_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_4_ccff_tail),
		.mem_out(mem_out[52:56]),
		.mem_outb(mem_outb[52:56]));

	cb_mux_size26_mem mem_top_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_5_ccff_tail),
		.mem_out(mem_out[57:61]),
		.mem_outb(mem_outb[57:61]));

	cb_mux_size26_mem mem_top_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_6_ccff_tail),
		.mem_out(mem_out[62:66]),
		.mem_outb(mem_outb[62:66]));

	cb_mux_size26_mem mem_top_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_7_ccff_tail),
		.mem_out(mem_out[67:71]),
		.mem_outb(mem_outb[67:71]));

	cb_mux_size26_mem mem_top_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_8_ccff_tail),
		.mem_out(mem_out[72:76]),
		.mem_outb(mem_outb[72:76]));

	cb_mux_size26_mem mem_top_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_9_ccff_tail),
		.mem_out(mem_out[77:81]),
		.mem_outb(mem_outb[77:81]));

	cb_mux_size26_mem mem_top_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_10_ccff_tail),
		.mem_out(mem_out[82:86]),
		.mem_outb(mem_outb[82:86]));

	cb_mux_size26_mem mem_top_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_11_ccff_tail),
		.mem_out(mem_out[87:91]),
		.mem_outb(mem_outb[87:91]));

	cb_mux_size26_mem mem_top_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_12_ccff_tail),
		.mem_out(mem_out[92:96]),
		.mem_outb(mem_outb[92:96]));

	cb_mux_size26_mem mem_top_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_13_ccff_tail),
		.mem_out(mem_out[97:101]),
		.mem_outb(mem_outb[97:101]));

	cb_mux_size26_mem mem_top_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_14_ccff_tail),
		.mem_out(mem_out[102:106]),
		.mem_outb(mem_outb[102:106]));

	cb_mux_size26_mem mem_top_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_15_ccff_tail),
		.mem_out(mem_out[107:111]),
		.mem_outb(mem_outb[107:111]));

	cb_mux_size26_mem mem_top_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_16_ccff_tail),
		.mem_out(mem_out[112:116]),
		.mem_outb(mem_outb[112:116]));

	cb_mux_size26_mem mem_top_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_17_ccff_tail),
		.mem_out(mem_out[117:121]),
		.mem_outb(mem_outb[117:121]));

	cb_mux_size26_mem mem_top_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_18_ccff_tail),
		.mem_out(mem_out[122:126]),
		.mem_outb(mem_outb[122:126]));

	cb_mux_size26_mem mem_top_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_19_ccff_tail),
		.mem_out(mem_out[127:131]),
		.mem_outb(mem_outb[127:131]));

	cb_mux_size26_mem mem_top_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_20_ccff_tail),
		.mem_out(mem_out[132:136]),
		.mem_outb(mem_outb[132:136]));

	cb_mux_size26_mem mem_top_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_21_ccff_tail),
		.mem_out(mem_out[137:141]),
		.mem_outb(mem_outb[137:141]));

	cb_mux_size26_mem mem_top_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_22_ccff_tail),
		.mem_out(mem_out[142:146]),
		.mem_outb(mem_outb[142:146]));

	cb_mux_size26_mem mem_top_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_23_ccff_tail),
		.mem_out(mem_out[147:151]),
		.mem_outb(mem_outb[147:151]));

	cb_mux_size26_mem mem_top_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_24_ccff_tail),
		.mem_out(mem_out[152:156]),
		.mem_outb(mem_outb[152:156]));

	cb_mux_size26_mem mem_top_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_25_ccff_tail),
		.mem_out(mem_out[157:161]),
		.mem_outb(mem_outb[157:161]));

	cb_mux_size26_mem mem_top_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_26_ccff_tail),
		.mem_out(mem_out[162:166]),
		.mem_outb(mem_outb[162:166]));

	cb_mux_size26_mem mem_top_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_27_ccff_tail),
		.mem_out(mem_out[167:171]),
		.mem_outb(mem_outb[167:171]));

	cb_mux_size26_mem mem_top_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_28_ccff_tail),
		.mem_out(mem_out[172:176]),
		.mem_outb(mem_outb[172:176]));

	cb_mux_size26_mem mem_top_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_29_ccff_tail),
		.mem_out(mem_out[177:181]),
		.mem_outb(mem_outb[177:181]));

endmodule
// ----- END Verilog module for cbx_4__config_group_mem_size206 -----




// ----- Verilog module for cbx_5__config_group_mem_size174 -----
module cbx_5__config_group_mem_size174(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:173] mem_out;
//----- OUTPUT PORTS -----
output [0:173] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size26_mem mem_top_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size26_mem_0_ccff_tail),
		.mem_out(mem_out[0:4]),
		.mem_outb(mem_outb[0:4]));

	cb_mux_size26_mem mem_top_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_1_ccff_tail),
		.mem_out(mem_out[5:9]),
		.mem_outb(mem_outb[5:9]));

	cb_mux_size26_mem mem_top_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_2_ccff_tail),
		.mem_out(mem_out[10:14]),
		.mem_outb(mem_outb[10:14]));

	cb_mux_size26_mem mem_top_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_3_ccff_tail),
		.mem_out(mem_out[15:19]),
		.mem_outb(mem_outb[15:19]));

	cb_mux_size26_mem mem_top_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_4_ccff_tail),
		.mem_out(mem_out[20:24]),
		.mem_outb(mem_outb[20:24]));

	cb_mux_size26_mem mem_top_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_5_ccff_tail),
		.mem_out(mem_out[25:29]),
		.mem_outb(mem_outb[25:29]));

	cb_mux_size26_mem mem_top_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_6_ccff_tail),
		.mem_out(mem_out[30:34]),
		.mem_outb(mem_outb[30:34]));

	cb_mux_size26_mem mem_top_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_7_ccff_tail),
		.mem_out(mem_out[35:39]),
		.mem_outb(mem_outb[35:39]));

	cb_mux_size26_mem mem_top_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_8_ccff_tail),
		.mem_out(mem_out[40:44]),
		.mem_outb(mem_outb[40:44]));

	cb_mux_size26_mem mem_top_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_9_ccff_tail),
		.mem_out(mem_out[45:49]),
		.mem_outb(mem_outb[45:49]));

	cb_mux_size26_mem mem_top_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_10_ccff_tail),
		.mem_out(mem_out[50:54]),
		.mem_outb(mem_outb[50:54]));

	cb_mux_size26_mem mem_top_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_11_ccff_tail),
		.mem_out(mem_out[55:59]),
		.mem_outb(mem_outb[55:59]));

	cb_mux_size26_mem mem_top_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_12_ccff_tail),
		.mem_out(mem_out[60:64]),
		.mem_outb(mem_outb[60:64]));

	cb_mux_size26_mem mem_top_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_13_ccff_tail),
		.mem_out(mem_out[65:69]),
		.mem_outb(mem_outb[65:69]));

	cb_mux_size26_mem mem_top_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_14_ccff_tail),
		.mem_out(mem_out[70:74]),
		.mem_outb(mem_outb[70:74]));

	cb_mux_size26_mem mem_top_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_15_ccff_tail),
		.mem_out(mem_out[75:79]),
		.mem_outb(mem_outb[75:79]));

	cb_mux_size26_mem mem_top_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_16_ccff_tail),
		.mem_out(mem_out[80:84]),
		.mem_outb(mem_outb[80:84]));

	cb_mux_size26_mem mem_top_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_17_ccff_tail),
		.mem_out(mem_out[85:89]),
		.mem_outb(mem_outb[85:89]));

	cb_mux_size26_mem mem_top_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_18_ccff_tail),
		.mem_out(mem_out[90:94]),
		.mem_outb(mem_outb[90:94]));

	cb_mux_size26_mem mem_top_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_19_ccff_tail),
		.mem_out(mem_out[95:99]),
		.mem_outb(mem_outb[95:99]));

	cb_mux_size26_mem mem_top_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_20_ccff_tail),
		.mem_out(mem_out[100:104]),
		.mem_outb(mem_outb[100:104]));

	cb_mux_size26_mem mem_top_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_21_ccff_tail),
		.mem_out(mem_out[105:109]),
		.mem_outb(mem_outb[105:109]));

	cb_mux_size26_mem mem_top_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_22_ccff_tail),
		.mem_out(mem_out[110:114]),
		.mem_outb(mem_outb[110:114]));

	cb_mux_size26_mem mem_top_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_23_ccff_tail),
		.mem_out(mem_out[115:119]),
		.mem_outb(mem_outb[115:119]));

	cb_mux_size26_mem mem_top_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_24_ccff_tail),
		.mem_out(mem_out[120:124]),
		.mem_outb(mem_outb[120:124]));

	cb_mux_size26_mem mem_top_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_25_ccff_tail),
		.mem_out(mem_out[125:129]),
		.mem_outb(mem_outb[125:129]));

	cb_mux_size26_mem mem_top_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_26_ccff_tail),
		.mem_out(mem_out[130:134]),
		.mem_outb(mem_outb[130:134]));

	cb_mux_size26_mem mem_top_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_27_ccff_tail),
		.mem_out(mem_out[135:139]),
		.mem_outb(mem_outb[135:139]));

	cb_mux_size26_mem mem_top_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_28_ccff_tail),
		.mem_out(mem_out[140:144]),
		.mem_outb(mem_outb[140:144]));

	cb_mux_size26_mem mem_top_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_29_ccff_tail),
		.mem_out(mem_out[145:149]),
		.mem_outb(mem_outb[145:149]));

	cb_mux_size8_mem mem_top_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[150:153]),
		.mem_outb(mem_outb[150:153]));

	cb_mux_size8_mem mem_top_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[154:157]),
		.mem_outb(mem_outb[154:157]));

	cb_mux_size8_mem mem_top_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[158:161]),
		.mem_outb(mem_outb[158:161]));

	cb_mux_size8_mem mem_top_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[162:165]),
		.mem_outb(mem_outb[162:165]));

	cb_mux_size8_mem mem_top_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[166:169]),
		.mem_outb(mem_outb[166:169]));

	cb_mux_size8_mem mem_top_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[170:173]),
		.mem_outb(mem_outb[170:173]));

endmodule
// ----- END Verilog module for cbx_5__config_group_mem_size174 -----




// ----- Verilog module for cbx_6__config_group_mem_size206 -----
module cbx_6__config_group_mem_size206(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:205] mem_out;
//----- OUTPUT PORTS -----
output [0:205] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size8_mem mem_bottom_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[0:3]),
		.mem_outb(mem_outb[0:3]));

	cb_mux_size8_mem mem_bottom_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[4:7]),
		.mem_outb(mem_outb[4:7]));

	cb_mux_size8_mem mem_bottom_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[8:11]),
		.mem_outb(mem_outb[8:11]));

	cb_mux_size8_mem mem_bottom_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[12:15]),
		.mem_outb(mem_outb[12:15]));

	cb_mux_size8_mem mem_bottom_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[16:19]),
		.mem_outb(mem_outb[16:19]));

	cb_mux_size8_mem mem_bottom_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[20:23]),
		.mem_outb(mem_outb[20:23]));

	cb_mux_size8_mem mem_bottom_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[24:27]),
		.mem_outb(mem_outb[24:27]));

	cb_mux_size8_mem mem_bottom_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[28:31]),
		.mem_outb(mem_outb[28:31]));

	cb_mux_size8_mem mem_top_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[182:185]),
		.mem_outb(mem_outb[182:185]));

	cb_mux_size8_mem mem_top_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[186:189]),
		.mem_outb(mem_outb[186:189]));

	cb_mux_size8_mem mem_top_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_10_ccff_tail),
		.mem_out(mem_out[190:193]),
		.mem_outb(mem_outb[190:193]));

	cb_mux_size8_mem mem_top_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_11_ccff_tail),
		.mem_out(mem_out[194:197]),
		.mem_outb(mem_outb[194:197]));

	cb_mux_size8_mem mem_top_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_12_ccff_tail),
		.mem_out(mem_out[198:201]),
		.mem_outb(mem_outb[198:201]));

	cb_mux_size8_mem mem_top_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_12_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[202:205]),
		.mem_outb(mem_outb[202:205]));

	cb_mux_size26_mem mem_top_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_0_ccff_tail),
		.mem_out(mem_out[32:36]),
		.mem_outb(mem_outb[32:36]));

	cb_mux_size26_mem mem_top_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_1_ccff_tail),
		.mem_out(mem_out[37:41]),
		.mem_outb(mem_outb[37:41]));

	cb_mux_size26_mem mem_top_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_2_ccff_tail),
		.mem_out(mem_out[42:46]),
		.mem_outb(mem_outb[42:46]));

	cb_mux_size26_mem mem_top_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_3_ccff_tail),
		.mem_out(mem_out[47:51]),
		.mem_outb(mem_outb[47:51]));

	cb_mux_size26_mem mem_top_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_4_ccff_tail),
		.mem_out(mem_out[52:56]),
		.mem_outb(mem_outb[52:56]));

	cb_mux_size26_mem mem_top_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_5_ccff_tail),
		.mem_out(mem_out[57:61]),
		.mem_outb(mem_outb[57:61]));

	cb_mux_size26_mem mem_top_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_6_ccff_tail),
		.mem_out(mem_out[62:66]),
		.mem_outb(mem_outb[62:66]));

	cb_mux_size26_mem mem_top_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_7_ccff_tail),
		.mem_out(mem_out[67:71]),
		.mem_outb(mem_outb[67:71]));

	cb_mux_size26_mem mem_top_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_8_ccff_tail),
		.mem_out(mem_out[72:76]),
		.mem_outb(mem_outb[72:76]));

	cb_mux_size26_mem mem_top_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_9_ccff_tail),
		.mem_out(mem_out[77:81]),
		.mem_outb(mem_outb[77:81]));

	cb_mux_size26_mem mem_top_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_10_ccff_tail),
		.mem_out(mem_out[82:86]),
		.mem_outb(mem_outb[82:86]));

	cb_mux_size26_mem mem_top_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_11_ccff_tail),
		.mem_out(mem_out[87:91]),
		.mem_outb(mem_outb[87:91]));

	cb_mux_size26_mem mem_top_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_12_ccff_tail),
		.mem_out(mem_out[92:96]),
		.mem_outb(mem_outb[92:96]));

	cb_mux_size26_mem mem_top_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_13_ccff_tail),
		.mem_out(mem_out[97:101]),
		.mem_outb(mem_outb[97:101]));

	cb_mux_size26_mem mem_top_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_14_ccff_tail),
		.mem_out(mem_out[102:106]),
		.mem_outb(mem_outb[102:106]));

	cb_mux_size26_mem mem_top_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_15_ccff_tail),
		.mem_out(mem_out[107:111]),
		.mem_outb(mem_outb[107:111]));

	cb_mux_size26_mem mem_top_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_16_ccff_tail),
		.mem_out(mem_out[112:116]),
		.mem_outb(mem_outb[112:116]));

	cb_mux_size26_mem mem_top_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_17_ccff_tail),
		.mem_out(mem_out[117:121]),
		.mem_outb(mem_outb[117:121]));

	cb_mux_size26_mem mem_top_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_18_ccff_tail),
		.mem_out(mem_out[122:126]),
		.mem_outb(mem_outb[122:126]));

	cb_mux_size26_mem mem_top_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_19_ccff_tail),
		.mem_out(mem_out[127:131]),
		.mem_outb(mem_outb[127:131]));

	cb_mux_size26_mem mem_top_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_20_ccff_tail),
		.mem_out(mem_out[132:136]),
		.mem_outb(mem_outb[132:136]));

	cb_mux_size26_mem mem_top_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_21_ccff_tail),
		.mem_out(mem_out[137:141]),
		.mem_outb(mem_outb[137:141]));

	cb_mux_size26_mem mem_top_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_22_ccff_tail),
		.mem_out(mem_out[142:146]),
		.mem_outb(mem_outb[142:146]));

	cb_mux_size26_mem mem_top_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_23_ccff_tail),
		.mem_out(mem_out[147:151]),
		.mem_outb(mem_outb[147:151]));

	cb_mux_size26_mem mem_top_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_24_ccff_tail),
		.mem_out(mem_out[152:156]),
		.mem_outb(mem_outb[152:156]));

	cb_mux_size26_mem mem_top_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_25_ccff_tail),
		.mem_out(mem_out[157:161]),
		.mem_outb(mem_outb[157:161]));

	cb_mux_size26_mem mem_top_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_26_ccff_tail),
		.mem_out(mem_out[162:166]),
		.mem_outb(mem_outb[162:166]));

	cb_mux_size26_mem mem_top_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_27_ccff_tail),
		.mem_out(mem_out[167:171]),
		.mem_outb(mem_outb[167:171]));

	cb_mux_size26_mem mem_top_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_28_ccff_tail),
		.mem_out(mem_out[172:176]),
		.mem_outb(mem_outb[172:176]));

	cb_mux_size26_mem mem_top_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size26_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size26_mem_29_ccff_tail),
		.mem_out(mem_out[177:181]),
		.mem_outb(mem_outb[177:181]));

endmodule
// ----- END Verilog module for cbx_6__config_group_mem_size206 -----




// ----- Verilog module for cby_1__config_group_mem_size224 -----
module cby_1__config_group_mem_size224(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:223] mem_out;
//----- OUTPUT PORTS -----
output [0:223] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size48_mem mem_right_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size48_mem_0_ccff_tail),
		.mem_out(mem_out[0:5]),
		.mem_outb(mem_outb[0:5]));

	cb_mux_size48_mem mem_right_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_1_ccff_tail),
		.mem_out(mem_out[11:16]),
		.mem_outb(mem_outb[11:16]));

	cb_mux_size48_mem mem_right_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_2_ccff_tail),
		.mem_out(mem_out[22:27]),
		.mem_outb(mem_outb[22:27]));

	cb_mux_size48_mem mem_right_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_3_ccff_tail),
		.mem_out(mem_out[33:38]),
		.mem_outb(mem_outb[33:38]));

	cb_mux_size48_mem mem_right_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_4_ccff_tail),
		.mem_out(mem_out[44:49]),
		.mem_outb(mem_outb[44:49]));

	cb_mux_size48_mem mem_right_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_5_ccff_tail),
		.mem_out(mem_out[55:60]),
		.mem_outb(mem_outb[55:60]));

	cb_mux_size48_mem mem_right_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_6_ccff_tail),
		.mem_out(mem_out[66:71]),
		.mem_outb(mem_outb[66:71]));

	cb_mux_size48_mem mem_right_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_7_ccff_tail),
		.mem_out(mem_out[77:82]),
		.mem_outb(mem_outb[77:82]));

	cb_mux_size48_mem mem_right_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_8_ccff_tail),
		.mem_out(mem_out[94:99]),
		.mem_outb(mem_outb[94:99]));

	cb_mux_size48_mem mem_right_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_9_ccff_tail),
		.mem_out(mem_out[111:116]),
		.mem_outb(mem_outb[111:116]));

	cb_mux_size48_mem mem_right_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_10_ccff_tail),
		.mem_out(mem_out[128:133]),
		.mem_outb(mem_outb[128:133]));

	cb_mux_size48_mem mem_right_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_11_ccff_tail),
		.mem_out(mem_out[145:150]),
		.mem_outb(mem_outb[145:150]));

	cb_mux_size48_mem mem_right_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_12_ccff_tail),
		.mem_out(mem_out[162:167]),
		.mem_outb(mem_outb[162:167]));

	cb_mux_size48_mem mem_right_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_13_ccff_tail),
		.mem_out(mem_out[179:184]),
		.mem_outb(mem_outb[179:184]));

	cb_mux_size48_mem mem_right_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_14_ccff_tail),
		.mem_out(mem_out[196:201]),
		.mem_outb(mem_outb[196:201]));

	cb_mux_size48_mem mem_right_ipin_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_15_ccff_tail),
		.mem_out(mem_out[213:218]),
		.mem_outb(mem_outb[213:218]));

	cb_mux_size16_mem mem_right_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_0_ccff_tail),
		.mem_out(mem_out[6:10]),
		.mem_outb(mem_outb[6:10]));

	cb_mux_size16_mem mem_right_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_1_ccff_tail),
		.mem_out(mem_out[17:21]),
		.mem_outb(mem_outb[17:21]));

	cb_mux_size16_mem mem_right_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_2_ccff_tail),
		.mem_out(mem_out[28:32]),
		.mem_outb(mem_outb[28:32]));

	cb_mux_size16_mem mem_right_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_3_ccff_tail),
		.mem_out(mem_out[39:43]),
		.mem_outb(mem_outb[39:43]));

	cb_mux_size16_mem mem_right_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_4_ccff_tail),
		.mem_out(mem_out[50:54]),
		.mem_outb(mem_outb[50:54]));

	cb_mux_size16_mem mem_right_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_5_ccff_tail),
		.mem_out(mem_out[61:65]),
		.mem_outb(mem_outb[61:65]));

	cb_mux_size16_mem mem_right_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_6_ccff_tail),
		.mem_out(mem_out[72:76]),
		.mem_outb(mem_outb[72:76]));

	cb_mux_size16_mem mem_right_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_7_ccff_tail),
		.mem_out(mem_out[83:87]),
		.mem_outb(mem_outb[83:87]));

	cb_mux_size16_mem mem_right_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_8_ccff_tail),
		.mem_out(mem_out[100:104]),
		.mem_outb(mem_outb[100:104]));

	cb_mux_size16_mem mem_right_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_9_ccff_tail),
		.mem_out(mem_out[117:121]),
		.mem_outb(mem_outb[117:121]));

	cb_mux_size16_mem mem_right_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_10_ccff_tail),
		.mem_out(mem_out[134:138]),
		.mem_outb(mem_outb[134:138]));

	cb_mux_size16_mem mem_right_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_11_ccff_tail),
		.mem_out(mem_out[151:155]),
		.mem_outb(mem_outb[151:155]));

	cb_mux_size16_mem mem_right_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_12_ccff_tail),
		.mem_out(mem_out[168:172]),
		.mem_outb(mem_outb[168:172]));

	cb_mux_size16_mem mem_right_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_13_ccff_tail),
		.mem_out(mem_out[185:189]),
		.mem_outb(mem_outb[185:189]));

	cb_mux_size16_mem mem_right_ipin_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_14_ccff_tail),
		.mem_out(mem_out[202:206]),
		.mem_outb(mem_outb[202:206]));

	cb_mux_size16_mem mem_right_ipin_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_15_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[219:223]),
		.mem_outb(mem_outb[219:223]));

	cb_mux_size56_mem mem_right_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_0_ccff_tail),
		.mem_out(mem_out[88:93]),
		.mem_outb(mem_outb[88:93]));

	cb_mux_size56_mem mem_right_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_1_ccff_tail),
		.mem_out(mem_out[105:110]),
		.mem_outb(mem_outb[105:110]));

	cb_mux_size56_mem mem_right_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_2_ccff_tail),
		.mem_out(mem_out[122:127]),
		.mem_outb(mem_outb[122:127]));

	cb_mux_size56_mem mem_right_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_3_ccff_tail),
		.mem_out(mem_out[139:144]),
		.mem_outb(mem_outb[139:144]));

	cb_mux_size56_mem mem_right_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_4_ccff_tail),
		.mem_out(mem_out[156:161]),
		.mem_outb(mem_outb[156:161]));

	cb_mux_size56_mem mem_right_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_5_ccff_tail),
		.mem_out(mem_out[173:178]),
		.mem_outb(mem_outb[173:178]));

	cb_mux_size56_mem mem_right_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_6_ccff_tail),
		.mem_out(mem_out[190:195]),
		.mem_outb(mem_outb[190:195]));

	cb_mux_size56_mem mem_right_ipin_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_7_ccff_tail),
		.mem_out(mem_out[207:212]),
		.mem_outb(mem_outb[207:212]));

endmodule
// ----- END Verilog module for cby_1__config_group_mem_size224 -----




// ----- Verilog module for cby_2__config_group_mem_size176 -----
module cby_2__config_group_mem_size176(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:175] mem_out;
//----- OUTPUT PORTS -----
output [0:175] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size48_mem mem_right_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size48_mem_0_ccff_tail),
		.mem_out(mem_out[0:5]),
		.mem_outb(mem_outb[0:5]));

	cb_mux_size48_mem mem_right_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_1_ccff_tail),
		.mem_out(mem_out[11:16]),
		.mem_outb(mem_outb[11:16]));

	cb_mux_size48_mem mem_right_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_2_ccff_tail),
		.mem_out(mem_out[22:27]),
		.mem_outb(mem_outb[22:27]));

	cb_mux_size48_mem mem_right_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_3_ccff_tail),
		.mem_out(mem_out[33:38]),
		.mem_outb(mem_outb[33:38]));

	cb_mux_size48_mem mem_right_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_4_ccff_tail),
		.mem_out(mem_out[44:49]),
		.mem_outb(mem_outb[44:49]));

	cb_mux_size48_mem mem_right_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_5_ccff_tail),
		.mem_out(mem_out[55:60]),
		.mem_outb(mem_outb[55:60]));

	cb_mux_size48_mem mem_right_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_6_ccff_tail),
		.mem_out(mem_out[66:71]),
		.mem_outb(mem_outb[66:71]));

	cb_mux_size48_mem mem_right_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_7_ccff_tail),
		.mem_out(mem_out[77:82]),
		.mem_outb(mem_outb[77:82]));

	cb_mux_size48_mem mem_right_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_8_ccff_tail),
		.mem_out(mem_out[88:93]),
		.mem_outb(mem_outb[88:93]));

	cb_mux_size48_mem mem_right_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_9_ccff_tail),
		.mem_out(mem_out[99:104]),
		.mem_outb(mem_outb[99:104]));

	cb_mux_size48_mem mem_right_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_10_ccff_tail),
		.mem_out(mem_out[110:115]),
		.mem_outb(mem_outb[110:115]));

	cb_mux_size48_mem mem_right_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_11_ccff_tail),
		.mem_out(mem_out[121:126]),
		.mem_outb(mem_outb[121:126]));

	cb_mux_size48_mem mem_right_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_12_ccff_tail),
		.mem_out(mem_out[132:137]),
		.mem_outb(mem_outb[132:137]));

	cb_mux_size48_mem mem_right_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_13_ccff_tail),
		.mem_out(mem_out[143:148]),
		.mem_outb(mem_outb[143:148]));

	cb_mux_size48_mem mem_right_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_14_ccff_tail),
		.mem_out(mem_out[154:159]),
		.mem_outb(mem_outb[154:159]));

	cb_mux_size48_mem mem_right_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_15_ccff_tail),
		.mem_out(mem_out[165:170]),
		.mem_outb(mem_outb[165:170]));

	cb_mux_size16_mem mem_right_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_0_ccff_tail),
		.mem_out(mem_out[6:10]),
		.mem_outb(mem_outb[6:10]));

	cb_mux_size16_mem mem_right_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_1_ccff_tail),
		.mem_out(mem_out[17:21]),
		.mem_outb(mem_outb[17:21]));

	cb_mux_size16_mem mem_right_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_2_ccff_tail),
		.mem_out(mem_out[28:32]),
		.mem_outb(mem_outb[28:32]));

	cb_mux_size16_mem mem_right_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_3_ccff_tail),
		.mem_out(mem_out[39:43]),
		.mem_outb(mem_outb[39:43]));

	cb_mux_size16_mem mem_right_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_4_ccff_tail),
		.mem_out(mem_out[50:54]),
		.mem_outb(mem_outb[50:54]));

	cb_mux_size16_mem mem_right_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_5_ccff_tail),
		.mem_out(mem_out[61:65]),
		.mem_outb(mem_outb[61:65]));

	cb_mux_size16_mem mem_right_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_6_ccff_tail),
		.mem_out(mem_out[72:76]),
		.mem_outb(mem_outb[72:76]));

	cb_mux_size16_mem mem_right_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_7_ccff_tail),
		.mem_out(mem_out[83:87]),
		.mem_outb(mem_outb[83:87]));

	cb_mux_size16_mem mem_right_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_8_ccff_tail),
		.mem_out(mem_out[94:98]),
		.mem_outb(mem_outb[94:98]));

	cb_mux_size16_mem mem_right_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_9_ccff_tail),
		.mem_out(mem_out[105:109]),
		.mem_outb(mem_outb[105:109]));

	cb_mux_size16_mem mem_right_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_10_ccff_tail),
		.mem_out(mem_out[116:120]),
		.mem_outb(mem_outb[116:120]));

	cb_mux_size16_mem mem_right_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_11_ccff_tail),
		.mem_out(mem_out[127:131]),
		.mem_outb(mem_outb[127:131]));

	cb_mux_size16_mem mem_right_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_12_ccff_tail),
		.mem_out(mem_out[138:142]),
		.mem_outb(mem_outb[138:142]));

	cb_mux_size16_mem mem_right_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_13_ccff_tail),
		.mem_out(mem_out[149:153]),
		.mem_outb(mem_outb[149:153]));

	cb_mux_size16_mem mem_right_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_14_ccff_tail),
		.mem_out(mem_out[160:164]),
		.mem_outb(mem_outb[160:164]));

	cb_mux_size16_mem mem_right_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_15_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[171:175]),
		.mem_outb(mem_outb[171:175]));

endmodule
// ----- END Verilog module for cby_2__config_group_mem_size176 -----




// ----- Verilog module for cby_3__config_group_mem_size336 -----
module cby_3__config_group_mem_size336(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:335] mem_out;
//----- OUTPUT PORTS -----
output [0:335] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size76_mem mem_right_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size76_mem_0_ccff_tail),
		.mem_out(mem_out[0:6]),
		.mem_outb(mem_outb[0:6]));

	cb_mux_size76_mem mem_right_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_1_ccff_tail),
		.mem_out(mem_out[7:13]),
		.mem_outb(mem_outb[7:13]));

	cb_mux_size76_mem mem_right_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_2_ccff_tail),
		.mem_out(mem_out[14:20]),
		.mem_outb(mem_outb[14:20]));

	cb_mux_size76_mem mem_right_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_3_ccff_tail),
		.mem_out(mem_out[21:27]),
		.mem_outb(mem_outb[21:27]));

	cb_mux_size76_mem mem_right_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_4_ccff_tail),
		.mem_out(mem_out[28:34]),
		.mem_outb(mem_outb[28:34]));

	cb_mux_size76_mem mem_right_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_5_ccff_tail),
		.mem_out(mem_out[35:41]),
		.mem_outb(mem_outb[35:41]));

	cb_mux_size76_mem mem_right_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_6_ccff_tail),
		.mem_out(mem_out[42:48]),
		.mem_outb(mem_outb[42:48]));

	cb_mux_size76_mem mem_right_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_7_ccff_tail),
		.mem_out(mem_out[49:55]),
		.mem_outb(mem_outb[49:55]));

	cb_mux_size76_mem mem_right_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_8_ccff_tail),
		.mem_out(mem_out[56:62]),
		.mem_outb(mem_outb[56:62]));

	cb_mux_size76_mem mem_right_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_9_ccff_tail),
		.mem_out(mem_out[63:69]),
		.mem_outb(mem_outb[63:69]));

	cb_mux_size76_mem mem_right_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_10_ccff_tail),
		.mem_out(mem_out[70:76]),
		.mem_outb(mem_outb[70:76]));

	cb_mux_size76_mem mem_right_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_11_ccff_tail),
		.mem_out(mem_out[77:83]),
		.mem_outb(mem_outb[77:83]));

	cb_mux_size76_mem mem_right_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_12_ccff_tail),
		.mem_out(mem_out[84:90]),
		.mem_outb(mem_outb[84:90]));

	cb_mux_size76_mem mem_right_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_13_ccff_tail),
		.mem_out(mem_out[91:97]),
		.mem_outb(mem_outb[91:97]));

	cb_mux_size76_mem mem_right_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_14_ccff_tail),
		.mem_out(mem_out[98:104]),
		.mem_outb(mem_outb[98:104]));

	cb_mux_size76_mem mem_right_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_15_ccff_tail),
		.mem_out(mem_out[105:111]),
		.mem_outb(mem_outb[105:111]));

	cb_mux_size76_mem mem_right_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_16_ccff_tail),
		.mem_out(mem_out[112:118]),
		.mem_outb(mem_outb[112:118]));

	cb_mux_size76_mem mem_right_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_17_ccff_tail),
		.mem_out(mem_out[119:125]),
		.mem_outb(mem_outb[119:125]));

	cb_mux_size76_mem mem_right_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_18_ccff_tail),
		.mem_out(mem_out[126:132]),
		.mem_outb(mem_outb[126:132]));

	cb_mux_size76_mem mem_right_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_19_ccff_tail),
		.mem_out(mem_out[133:139]),
		.mem_outb(mem_outb[133:139]));

	cb_mux_size76_mem mem_right_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_20_ccff_tail),
		.mem_out(mem_out[140:146]),
		.mem_outb(mem_outb[140:146]));

	cb_mux_size76_mem mem_right_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_21_ccff_tail),
		.mem_out(mem_out[147:153]),
		.mem_outb(mem_outb[147:153]));

	cb_mux_size76_mem mem_right_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_22_ccff_tail),
		.mem_out(mem_out[154:160]),
		.mem_outb(mem_outb[154:160]));

	cb_mux_size76_mem mem_right_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_23_ccff_tail),
		.mem_out(mem_out[161:167]),
		.mem_outb(mem_outb[161:167]));

	cb_mux_size76_mem mem_right_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_24_ccff_tail),
		.mem_out(mem_out[168:174]),
		.mem_outb(mem_outb[168:174]));

	cb_mux_size76_mem mem_right_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_25_ccff_tail),
		.mem_out(mem_out[175:181]),
		.mem_outb(mem_outb[175:181]));

	cb_mux_size76_mem mem_right_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_26_ccff_tail),
		.mem_out(mem_out[182:188]),
		.mem_outb(mem_outb[182:188]));

	cb_mux_size76_mem mem_right_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_27_ccff_tail),
		.mem_out(mem_out[189:195]),
		.mem_outb(mem_outb[189:195]));

	cb_mux_size76_mem mem_right_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_28_ccff_tail),
		.mem_out(mem_out[196:202]),
		.mem_outb(mem_outb[196:202]));

	cb_mux_size76_mem mem_right_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_29_ccff_tail),
		.mem_out(mem_out[203:209]),
		.mem_outb(mem_outb[203:209]));

	cb_mux_size48_mem mem_right_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_0_ccff_tail),
		.mem_out(mem_out[210:215]),
		.mem_outb(mem_outb[210:215]));

	cb_mux_size48_mem mem_right_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_1_ccff_tail),
		.mem_out(mem_out[221:226]),
		.mem_outb(mem_outb[221:226]));

	cb_mux_size48_mem mem_right_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_2_ccff_tail),
		.mem_out(mem_out[238:243]),
		.mem_outb(mem_outb[238:243]));

	cb_mux_size48_mem mem_right_ipin_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_3_ccff_tail),
		.mem_out(mem_out[255:260]),
		.mem_outb(mem_outb[255:260]));

	cb_mux_size16_mem mem_right_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_0_ccff_tail),
		.mem_out(mem_out[216:220]),
		.mem_outb(mem_outb[216:220]));

	cb_mux_size16_mem mem_right_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_1_ccff_tail),
		.mem_out(mem_out[233:237]),
		.mem_outb(mem_outb[233:237]));

	cb_mux_size16_mem mem_right_ipin_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_2_ccff_tail),
		.mem_out(mem_out[250:254]),
		.mem_outb(mem_outb[250:254]));

	cb_mux_size16_mem mem_right_ipin_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_3_ccff_tail),
		.mem_out(mem_out[267:271]),
		.mem_outb(mem_outb[267:271]));

	cb_mux_size56_mem mem_right_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_0_ccff_tail),
		.mem_out(mem_out[227:232]),
		.mem_outb(mem_outb[227:232]));

	cb_mux_size56_mem mem_right_ipin_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_1_ccff_tail),
		.mem_out(mem_out[244:249]),
		.mem_outb(mem_outb[244:249]));

	cb_mux_size56_mem mem_right_ipin_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_2_ccff_tail),
		.mem_out(mem_out[261:266]),
		.mem_outb(mem_outb[261:266]));

	cb_mux_size8_mem mem_right_ipin_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[272:275]),
		.mem_outb(mem_outb[272:275]));

	cb_mux_size8_mem mem_right_ipin_42 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[276:279]),
		.mem_outb(mem_outb[276:279]));

	cb_mux_size8_mem mem_right_ipin_43 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[280:283]),
		.mem_outb(mem_outb[280:283]));

	cb_mux_size8_mem mem_right_ipin_44 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[284:287]),
		.mem_outb(mem_outb[284:287]));

	cb_mux_size8_mem mem_right_ipin_45 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[288:291]),
		.mem_outb(mem_outb[288:291]));

	cb_mux_size8_mem mem_right_ipin_46 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[292:295]),
		.mem_outb(mem_outb[292:295]));

	cb_mux_size8_mem mem_right_ipin_47 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[296:299]),
		.mem_outb(mem_outb[296:299]));

	cb_mux_size8_mem mem_right_ipin_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[300:303]),
		.mem_outb(mem_outb[300:303]));

	cb_mux_size8_mem mem_right_ipin_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[304:307]),
		.mem_outb(mem_outb[304:307]));

	cb_mux_size8_mem mem_right_ipin_50 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[308:311]),
		.mem_outb(mem_outb[308:311]));

	cb_mux_size8_mem mem_right_ipin_51 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_10_ccff_tail),
		.mem_out(mem_out[312:315]),
		.mem_outb(mem_outb[312:315]));

	cb_mux_size8_mem mem_right_ipin_52 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_11_ccff_tail),
		.mem_out(mem_out[316:319]),
		.mem_outb(mem_outb[316:319]));

	cb_mux_size8_mem mem_right_ipin_53 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_12_ccff_tail),
		.mem_out(mem_out[320:323]),
		.mem_outb(mem_outb[320:323]));

	cb_mux_size8_mem mem_right_ipin_54 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_13_ccff_tail),
		.mem_out(mem_out[324:327]),
		.mem_outb(mem_outb[324:327]));

	cb_mux_size8_mem mem_right_ipin_55 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_14_ccff_tail),
		.mem_out(mem_out[328:331]),
		.mem_outb(mem_outb[328:331]));

	cb_mux_size8_mem mem_right_ipin_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_14_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[332:335]),
		.mem_outb(mem_outb[332:335]));

endmodule
// ----- END Verilog module for cby_3__config_group_mem_size336 -----




// ----- Verilog module for cby_4__config_group_mem_size336 -----
module cby_4__config_group_mem_size336(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:335] mem_out;
//----- OUTPUT PORTS -----
output [0:335] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size76_mem mem_right_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size76_mem_0_ccff_tail),
		.mem_out(mem_out[0:6]),
		.mem_outb(mem_outb[0:6]));

	cb_mux_size76_mem mem_right_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_1_ccff_tail),
		.mem_out(mem_out[7:13]),
		.mem_outb(mem_outb[7:13]));

	cb_mux_size76_mem mem_right_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_2_ccff_tail),
		.mem_out(mem_out[14:20]),
		.mem_outb(mem_outb[14:20]));

	cb_mux_size76_mem mem_right_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_3_ccff_tail),
		.mem_out(mem_out[21:27]),
		.mem_outb(mem_outb[21:27]));

	cb_mux_size76_mem mem_right_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_4_ccff_tail),
		.mem_out(mem_out[28:34]),
		.mem_outb(mem_outb[28:34]));

	cb_mux_size76_mem mem_right_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_5_ccff_tail),
		.mem_out(mem_out[35:41]),
		.mem_outb(mem_outb[35:41]));

	cb_mux_size76_mem mem_right_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_6_ccff_tail),
		.mem_out(mem_out[42:48]),
		.mem_outb(mem_outb[42:48]));

	cb_mux_size76_mem mem_right_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_7_ccff_tail),
		.mem_out(mem_out[49:55]),
		.mem_outb(mem_outb[49:55]));

	cb_mux_size76_mem mem_right_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_8_ccff_tail),
		.mem_out(mem_out[56:62]),
		.mem_outb(mem_outb[56:62]));

	cb_mux_size76_mem mem_right_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_9_ccff_tail),
		.mem_out(mem_out[63:69]),
		.mem_outb(mem_outb[63:69]));

	cb_mux_size76_mem mem_right_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_10_ccff_tail),
		.mem_out(mem_out[70:76]),
		.mem_outb(mem_outb[70:76]));

	cb_mux_size76_mem mem_right_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_11_ccff_tail),
		.mem_out(mem_out[77:83]),
		.mem_outb(mem_outb[77:83]));

	cb_mux_size76_mem mem_right_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_12_ccff_tail),
		.mem_out(mem_out[84:90]),
		.mem_outb(mem_outb[84:90]));

	cb_mux_size76_mem mem_right_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_13_ccff_tail),
		.mem_out(mem_out[91:97]),
		.mem_outb(mem_outb[91:97]));

	cb_mux_size76_mem mem_right_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_14_ccff_tail),
		.mem_out(mem_out[98:104]),
		.mem_outb(mem_outb[98:104]));

	cb_mux_size76_mem mem_right_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_15_ccff_tail),
		.mem_out(mem_out[105:111]),
		.mem_outb(mem_outb[105:111]));

	cb_mux_size76_mem mem_right_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_16_ccff_tail),
		.mem_out(mem_out[112:118]),
		.mem_outb(mem_outb[112:118]));

	cb_mux_size76_mem mem_right_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_17_ccff_tail),
		.mem_out(mem_out[119:125]),
		.mem_outb(mem_outb[119:125]));

	cb_mux_size76_mem mem_right_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_18_ccff_tail),
		.mem_out(mem_out[126:132]),
		.mem_outb(mem_outb[126:132]));

	cb_mux_size76_mem mem_right_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_19_ccff_tail),
		.mem_out(mem_out[133:139]),
		.mem_outb(mem_outb[133:139]));

	cb_mux_size76_mem mem_right_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_20_ccff_tail),
		.mem_out(mem_out[140:146]),
		.mem_outb(mem_outb[140:146]));

	cb_mux_size76_mem mem_right_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_21_ccff_tail),
		.mem_out(mem_out[147:153]),
		.mem_outb(mem_outb[147:153]));

	cb_mux_size76_mem mem_right_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_22_ccff_tail),
		.mem_out(mem_out[154:160]),
		.mem_outb(mem_outb[154:160]));

	cb_mux_size76_mem mem_right_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_23_ccff_tail),
		.mem_out(mem_out[161:167]),
		.mem_outb(mem_outb[161:167]));

	cb_mux_size76_mem mem_right_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_24_ccff_tail),
		.mem_out(mem_out[168:174]),
		.mem_outb(mem_outb[168:174]));

	cb_mux_size76_mem mem_right_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_25_ccff_tail),
		.mem_out(mem_out[175:181]),
		.mem_outb(mem_outb[175:181]));

	cb_mux_size76_mem mem_right_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_26_ccff_tail),
		.mem_out(mem_out[182:188]),
		.mem_outb(mem_outb[182:188]));

	cb_mux_size76_mem mem_right_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_27_ccff_tail),
		.mem_out(mem_out[189:195]),
		.mem_outb(mem_outb[189:195]));

	cb_mux_size76_mem mem_right_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_28_ccff_tail),
		.mem_out(mem_out[196:202]),
		.mem_outb(mem_outb[196:202]));

	cb_mux_size76_mem mem_right_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_29_ccff_tail),
		.mem_out(mem_out[203:209]),
		.mem_outb(mem_outb[203:209]));

	cb_mux_size48_mem mem_right_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_0_ccff_tail),
		.mem_out(mem_out[210:215]),
		.mem_outb(mem_outb[210:215]));

	cb_mux_size48_mem mem_right_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_1_ccff_tail),
		.mem_out(mem_out[221:226]),
		.mem_outb(mem_outb[221:226]));

	cb_mux_size48_mem mem_right_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_2_ccff_tail),
		.mem_out(mem_out[238:243]),
		.mem_outb(mem_outb[238:243]));

	cb_mux_size48_mem mem_right_ipin_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_3_ccff_tail),
		.mem_out(mem_out[255:260]),
		.mem_outb(mem_outb[255:260]));

	cb_mux_size16_mem mem_right_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_0_ccff_tail),
		.mem_out(mem_out[216:220]),
		.mem_outb(mem_outb[216:220]));

	cb_mux_size16_mem mem_right_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_1_ccff_tail),
		.mem_out(mem_out[233:237]),
		.mem_outb(mem_outb[233:237]));

	cb_mux_size16_mem mem_right_ipin_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_2_ccff_tail),
		.mem_out(mem_out[250:254]),
		.mem_outb(mem_outb[250:254]));

	cb_mux_size16_mem mem_right_ipin_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_3_ccff_tail),
		.mem_out(mem_out[267:271]),
		.mem_outb(mem_outb[267:271]));

	cb_mux_size56_mem mem_right_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_0_ccff_tail),
		.mem_out(mem_out[227:232]),
		.mem_outb(mem_outb[227:232]));

	cb_mux_size56_mem mem_right_ipin_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_1_ccff_tail),
		.mem_out(mem_out[244:249]),
		.mem_outb(mem_outb[244:249]));

	cb_mux_size56_mem mem_right_ipin_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_2_ccff_tail),
		.mem_out(mem_out[261:266]),
		.mem_outb(mem_outb[261:266]));

	cb_mux_size8_mem mem_right_ipin_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[272:275]),
		.mem_outb(mem_outb[272:275]));

	cb_mux_size8_mem mem_right_ipin_42 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[276:279]),
		.mem_outb(mem_outb[276:279]));

	cb_mux_size8_mem mem_right_ipin_43 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[280:283]),
		.mem_outb(mem_outb[280:283]));

	cb_mux_size8_mem mem_right_ipin_44 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[284:287]),
		.mem_outb(mem_outb[284:287]));

	cb_mux_size8_mem mem_right_ipin_45 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[288:291]),
		.mem_outb(mem_outb[288:291]));

	cb_mux_size8_mem mem_right_ipin_46 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[292:295]),
		.mem_outb(mem_outb[292:295]));

	cb_mux_size8_mem mem_right_ipin_47 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[296:299]),
		.mem_outb(mem_outb[296:299]));

	cb_mux_size8_mem mem_right_ipin_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[300:303]),
		.mem_outb(mem_outb[300:303]));

	cb_mux_size8_mem mem_right_ipin_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[304:307]),
		.mem_outb(mem_outb[304:307]));

	cb_mux_size8_mem mem_right_ipin_50 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[308:311]),
		.mem_outb(mem_outb[308:311]));

	cb_mux_size8_mem mem_right_ipin_51 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_10_ccff_tail),
		.mem_out(mem_out[312:315]),
		.mem_outb(mem_outb[312:315]));

	cb_mux_size8_mem mem_right_ipin_52 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_11_ccff_tail),
		.mem_out(mem_out[316:319]),
		.mem_outb(mem_outb[316:319]));

	cb_mux_size8_mem mem_right_ipin_53 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_12_ccff_tail),
		.mem_out(mem_out[320:323]),
		.mem_outb(mem_outb[320:323]));

	cb_mux_size8_mem mem_right_ipin_54 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_13_ccff_tail),
		.mem_out(mem_out[324:327]),
		.mem_outb(mem_outb[324:327]));

	cb_mux_size8_mem mem_right_ipin_55 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_14_ccff_tail),
		.mem_out(mem_out[328:331]),
		.mem_outb(mem_outb[328:331]));

	cb_mux_size8_mem mem_right_ipin_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_14_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[332:335]),
		.mem_outb(mem_outb[332:335]));

endmodule
// ----- END Verilog module for cby_4__config_group_mem_size336 -----




// ----- Verilog module for cby_5__config_group_mem_size560 -----
module cby_5__config_group_mem_size560(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:559] mem_out;
//----- OUTPUT PORTS -----
output [0:559] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size48_mem mem_left_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size48_mem_0_ccff_tail),
		.mem_out(mem_out[0:5]),
		.mem_outb(mem_outb[0:5]));

	cb_mux_size48_mem mem_left_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_1_ccff_tail),
		.mem_out(mem_out[11:16]),
		.mem_outb(mem_outb[11:16]));

	cb_mux_size48_mem mem_left_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_2_ccff_tail),
		.mem_out(mem_out[22:27]),
		.mem_outb(mem_outb[22:27]));

	cb_mux_size48_mem mem_left_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_3_ccff_tail),
		.mem_out(mem_out[33:38]),
		.mem_outb(mem_outb[33:38]));

	cb_mux_size48_mem mem_left_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_4_ccff_tail),
		.mem_out(mem_out[44:49]),
		.mem_outb(mem_outb[44:49]));

	cb_mux_size48_mem mem_left_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_5_ccff_tail),
		.mem_out(mem_out[55:60]),
		.mem_outb(mem_outb[55:60]));

	cb_mux_size48_mem mem_left_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_6_ccff_tail),
		.mem_out(mem_out[66:71]),
		.mem_outb(mem_outb[66:71]));

	cb_mux_size48_mem mem_left_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_7_ccff_tail),
		.mem_out(mem_out[77:82]),
		.mem_outb(mem_outb[77:82]));

	cb_mux_size48_mem mem_left_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_8_ccff_tail),
		.mem_out(mem_out[94:99]),
		.mem_outb(mem_outb[94:99]));

	cb_mux_size48_mem mem_left_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_9_ccff_tail),
		.mem_out(mem_out[111:116]),
		.mem_outb(mem_outb[111:116]));

	cb_mux_size48_mem mem_left_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_10_ccff_tail),
		.mem_out(mem_out[128:133]),
		.mem_outb(mem_outb[128:133]));

	cb_mux_size48_mem mem_left_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_11_ccff_tail),
		.mem_out(mem_out[145:150]),
		.mem_outb(mem_outb[145:150]));

	cb_mux_size48_mem mem_left_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_12_ccff_tail),
		.mem_out(mem_out[162:167]),
		.mem_outb(mem_outb[162:167]));

	cb_mux_size48_mem mem_left_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_13_ccff_tail),
		.mem_out(mem_out[179:184]),
		.mem_outb(mem_outb[179:184]));

	cb_mux_size48_mem mem_left_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_14_ccff_tail),
		.mem_out(mem_out[196:201]),
		.mem_outb(mem_outb[196:201]));

	cb_mux_size48_mem mem_left_ipin_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_15_ccff_tail),
		.mem_out(mem_out[213:218]),
		.mem_outb(mem_outb[213:218]));

	cb_mux_size48_mem mem_right_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_16_ccff_tail),
		.mem_out(mem_out[434:439]),
		.mem_outb(mem_outb[434:439]));

	cb_mux_size48_mem mem_right_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_17_ccff_tail),
		.mem_out(mem_out[445:450]),
		.mem_outb(mem_outb[445:450]));

	cb_mux_size48_mem mem_right_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_18_ccff_tail),
		.mem_out(mem_out[462:467]),
		.mem_outb(mem_outb[462:467]));

	cb_mux_size48_mem mem_right_ipin_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_19_ccff_tail),
		.mem_out(mem_out[479:484]),
		.mem_outb(mem_outb[479:484]));

	cb_mux_size16_mem mem_left_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_0_ccff_tail),
		.mem_out(mem_out[6:10]),
		.mem_outb(mem_outb[6:10]));

	cb_mux_size16_mem mem_left_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_1_ccff_tail),
		.mem_out(mem_out[17:21]),
		.mem_outb(mem_outb[17:21]));

	cb_mux_size16_mem mem_left_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_2_ccff_tail),
		.mem_out(mem_out[28:32]),
		.mem_outb(mem_outb[28:32]));

	cb_mux_size16_mem mem_left_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_3_ccff_tail),
		.mem_out(mem_out[39:43]),
		.mem_outb(mem_outb[39:43]));

	cb_mux_size16_mem mem_left_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_4_ccff_tail),
		.mem_out(mem_out[50:54]),
		.mem_outb(mem_outb[50:54]));

	cb_mux_size16_mem mem_left_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_5_ccff_tail),
		.mem_out(mem_out[61:65]),
		.mem_outb(mem_outb[61:65]));

	cb_mux_size16_mem mem_left_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_6_ccff_tail),
		.mem_out(mem_out[72:76]),
		.mem_outb(mem_outb[72:76]));

	cb_mux_size16_mem mem_left_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_7_ccff_tail),
		.mem_out(mem_out[83:87]),
		.mem_outb(mem_outb[83:87]));

	cb_mux_size16_mem mem_left_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_8_ccff_tail),
		.mem_out(mem_out[100:104]),
		.mem_outb(mem_outb[100:104]));

	cb_mux_size16_mem mem_left_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_9_ccff_tail),
		.mem_out(mem_out[117:121]),
		.mem_outb(mem_outb[117:121]));

	cb_mux_size16_mem mem_left_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_10_ccff_tail),
		.mem_out(mem_out[134:138]),
		.mem_outb(mem_outb[134:138]));

	cb_mux_size16_mem mem_left_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_11_ccff_tail),
		.mem_out(mem_out[151:155]),
		.mem_outb(mem_outb[151:155]));

	cb_mux_size16_mem mem_left_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_12_ccff_tail),
		.mem_out(mem_out[168:172]),
		.mem_outb(mem_outb[168:172]));

	cb_mux_size16_mem mem_left_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_13_ccff_tail),
		.mem_out(mem_out[185:189]),
		.mem_outb(mem_outb[185:189]));

	cb_mux_size16_mem mem_left_ipin_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_14_ccff_tail),
		.mem_out(mem_out[202:206]),
		.mem_outb(mem_outb[202:206]));

	cb_mux_size16_mem mem_left_ipin_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_15_ccff_tail),
		.mem_out(mem_out[219:223]),
		.mem_outb(mem_outb[219:223]));

	cb_mux_size16_mem mem_right_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_16_ccff_tail),
		.mem_out(mem_out[440:444]),
		.mem_outb(mem_outb[440:444]));

	cb_mux_size16_mem mem_right_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_17_ccff_tail),
		.mem_out(mem_out[457:461]),
		.mem_outb(mem_outb[457:461]));

	cb_mux_size16_mem mem_right_ipin_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_18_ccff_tail),
		.mem_out(mem_out[474:478]),
		.mem_outb(mem_outb[474:478]));

	cb_mux_size16_mem mem_right_ipin_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_19_ccff_tail),
		.mem_out(mem_out[491:495]),
		.mem_outb(mem_outb[491:495]));

	cb_mux_size56_mem mem_left_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_0_ccff_tail),
		.mem_out(mem_out[88:93]),
		.mem_outb(mem_outb[88:93]));

	cb_mux_size56_mem mem_left_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_1_ccff_tail),
		.mem_out(mem_out[105:110]),
		.mem_outb(mem_outb[105:110]));

	cb_mux_size56_mem mem_left_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_2_ccff_tail),
		.mem_out(mem_out[122:127]),
		.mem_outb(mem_outb[122:127]));

	cb_mux_size56_mem mem_left_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_3_ccff_tail),
		.mem_out(mem_out[139:144]),
		.mem_outb(mem_outb[139:144]));

	cb_mux_size56_mem mem_left_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_4_ccff_tail),
		.mem_out(mem_out[156:161]),
		.mem_outb(mem_outb[156:161]));

	cb_mux_size56_mem mem_left_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_5_ccff_tail),
		.mem_out(mem_out[173:178]),
		.mem_outb(mem_outb[173:178]));

	cb_mux_size56_mem mem_left_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_6_ccff_tail),
		.mem_out(mem_out[190:195]),
		.mem_outb(mem_outb[190:195]));

	cb_mux_size56_mem mem_left_ipin_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_7_ccff_tail),
		.mem_out(mem_out[207:212]),
		.mem_outb(mem_outb[207:212]));

	cb_mux_size56_mem mem_right_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_8_ccff_tail),
		.mem_out(mem_out[451:456]),
		.mem_outb(mem_outb[451:456]));

	cb_mux_size56_mem mem_right_ipin_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_9_ccff_tail),
		.mem_out(mem_out[468:473]),
		.mem_outb(mem_outb[468:473]));

	cb_mux_size56_mem mem_right_ipin_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_10_ccff_tail),
		.mem_out(mem_out[485:490]),
		.mem_outb(mem_outb[485:490]));

	cb_mux_size76_mem mem_right_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_0_ccff_tail),
		.mem_out(mem_out[224:230]),
		.mem_outb(mem_outb[224:230]));

	cb_mux_size76_mem mem_right_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_1_ccff_tail),
		.mem_out(mem_out[231:237]),
		.mem_outb(mem_outb[231:237]));

	cb_mux_size76_mem mem_right_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_2_ccff_tail),
		.mem_out(mem_out[238:244]),
		.mem_outb(mem_outb[238:244]));

	cb_mux_size76_mem mem_right_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_3_ccff_tail),
		.mem_out(mem_out[245:251]),
		.mem_outb(mem_outb[245:251]));

	cb_mux_size76_mem mem_right_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_4_ccff_tail),
		.mem_out(mem_out[252:258]),
		.mem_outb(mem_outb[252:258]));

	cb_mux_size76_mem mem_right_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_5_ccff_tail),
		.mem_out(mem_out[259:265]),
		.mem_outb(mem_outb[259:265]));

	cb_mux_size76_mem mem_right_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_6_ccff_tail),
		.mem_out(mem_out[266:272]),
		.mem_outb(mem_outb[266:272]));

	cb_mux_size76_mem mem_right_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_7_ccff_tail),
		.mem_out(mem_out[273:279]),
		.mem_outb(mem_outb[273:279]));

	cb_mux_size76_mem mem_right_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_8_ccff_tail),
		.mem_out(mem_out[280:286]),
		.mem_outb(mem_outb[280:286]));

	cb_mux_size76_mem mem_right_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_9_ccff_tail),
		.mem_out(mem_out[287:293]),
		.mem_outb(mem_outb[287:293]));

	cb_mux_size76_mem mem_right_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_10_ccff_tail),
		.mem_out(mem_out[294:300]),
		.mem_outb(mem_outb[294:300]));

	cb_mux_size76_mem mem_right_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_11_ccff_tail),
		.mem_out(mem_out[301:307]),
		.mem_outb(mem_outb[301:307]));

	cb_mux_size76_mem mem_right_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_12_ccff_tail),
		.mem_out(mem_out[308:314]),
		.mem_outb(mem_outb[308:314]));

	cb_mux_size76_mem mem_right_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_13_ccff_tail),
		.mem_out(mem_out[315:321]),
		.mem_outb(mem_outb[315:321]));

	cb_mux_size76_mem mem_right_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_14_ccff_tail),
		.mem_out(mem_out[322:328]),
		.mem_outb(mem_outb[322:328]));

	cb_mux_size76_mem mem_right_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_15_ccff_tail),
		.mem_out(mem_out[329:335]),
		.mem_outb(mem_outb[329:335]));

	cb_mux_size76_mem mem_right_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_16_ccff_tail),
		.mem_out(mem_out[336:342]),
		.mem_outb(mem_outb[336:342]));

	cb_mux_size76_mem mem_right_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_17_ccff_tail),
		.mem_out(mem_out[343:349]),
		.mem_outb(mem_outb[343:349]));

	cb_mux_size76_mem mem_right_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_18_ccff_tail),
		.mem_out(mem_out[350:356]),
		.mem_outb(mem_outb[350:356]));

	cb_mux_size76_mem mem_right_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_19_ccff_tail),
		.mem_out(mem_out[357:363]),
		.mem_outb(mem_outb[357:363]));

	cb_mux_size76_mem mem_right_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_20_ccff_tail),
		.mem_out(mem_out[364:370]),
		.mem_outb(mem_outb[364:370]));

	cb_mux_size76_mem mem_right_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_21_ccff_tail),
		.mem_out(mem_out[371:377]),
		.mem_outb(mem_outb[371:377]));

	cb_mux_size76_mem mem_right_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_22_ccff_tail),
		.mem_out(mem_out[378:384]),
		.mem_outb(mem_outb[378:384]));

	cb_mux_size76_mem mem_right_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_23_ccff_tail),
		.mem_out(mem_out[385:391]),
		.mem_outb(mem_outb[385:391]));

	cb_mux_size76_mem mem_right_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_24_ccff_tail),
		.mem_out(mem_out[392:398]),
		.mem_outb(mem_outb[392:398]));

	cb_mux_size76_mem mem_right_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_25_ccff_tail),
		.mem_out(mem_out[399:405]),
		.mem_outb(mem_outb[399:405]));

	cb_mux_size76_mem mem_right_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_26_ccff_tail),
		.mem_out(mem_out[406:412]),
		.mem_outb(mem_outb[406:412]));

	cb_mux_size76_mem mem_right_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_27_ccff_tail),
		.mem_out(mem_out[413:419]),
		.mem_outb(mem_outb[413:419]));

	cb_mux_size76_mem mem_right_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_28_ccff_tail),
		.mem_out(mem_out[420:426]),
		.mem_outb(mem_outb[420:426]));

	cb_mux_size76_mem mem_right_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_29_ccff_tail),
		.mem_out(mem_out[427:433]),
		.mem_outb(mem_outb[427:433]));

	cb_mux_size8_mem mem_right_ipin_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[496:499]),
		.mem_outb(mem_outb[496:499]));

	cb_mux_size8_mem mem_right_ipin_42 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[500:503]),
		.mem_outb(mem_outb[500:503]));

	cb_mux_size8_mem mem_right_ipin_43 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[504:507]),
		.mem_outb(mem_outb[504:507]));

	cb_mux_size8_mem mem_right_ipin_44 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[508:511]),
		.mem_outb(mem_outb[508:511]));

	cb_mux_size8_mem mem_right_ipin_45 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[512:515]),
		.mem_outb(mem_outb[512:515]));

	cb_mux_size8_mem mem_right_ipin_46 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[516:519]),
		.mem_outb(mem_outb[516:519]));

	cb_mux_size8_mem mem_right_ipin_47 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[520:523]),
		.mem_outb(mem_outb[520:523]));

	cb_mux_size8_mem mem_right_ipin_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[524:527]),
		.mem_outb(mem_outb[524:527]));

	cb_mux_size8_mem mem_right_ipin_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[528:531]),
		.mem_outb(mem_outb[528:531]));

	cb_mux_size8_mem mem_right_ipin_50 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[532:535]),
		.mem_outb(mem_outb[532:535]));

	cb_mux_size8_mem mem_right_ipin_51 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_10_ccff_tail),
		.mem_out(mem_out[536:539]),
		.mem_outb(mem_outb[536:539]));

	cb_mux_size8_mem mem_right_ipin_52 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_11_ccff_tail),
		.mem_out(mem_out[540:543]),
		.mem_outb(mem_outb[540:543]));

	cb_mux_size8_mem mem_right_ipin_53 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_12_ccff_tail),
		.mem_out(mem_out[544:547]),
		.mem_outb(mem_outb[544:547]));

	cb_mux_size8_mem mem_right_ipin_54 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_13_ccff_tail),
		.mem_out(mem_out[548:551]),
		.mem_outb(mem_outb[548:551]));

	cb_mux_size8_mem mem_right_ipin_55 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_14_ccff_tail),
		.mem_out(mem_out[552:555]),
		.mem_outb(mem_outb[552:555]));

	cb_mux_size8_mem mem_right_ipin_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_14_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[556:559]),
		.mem_outb(mem_outb[556:559]));

endmodule
// ----- END Verilog module for cby_5__config_group_mem_size560 -----




// ----- Verilog module for cby_6__config_group_mem_size560 -----
module cby_6__config_group_mem_size560(config_enable,
                                       prog_reset,
                                       prog_clk,
                                       ccff_head,
                                       mem_out,
                                       mem_outb,
                                       ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:559] mem_out;
//----- OUTPUT PORTS -----
output [0:559] mem_outb;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	cb_mux_size48_mem mem_left_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(cb_mux_size48_mem_0_ccff_tail),
		.mem_out(mem_out[0:5]),
		.mem_outb(mem_outb[0:5]));

	cb_mux_size48_mem mem_left_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_1_ccff_tail),
		.mem_out(mem_out[11:16]),
		.mem_outb(mem_outb[11:16]));

	cb_mux_size48_mem mem_left_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_2_ccff_tail),
		.mem_out(mem_out[22:27]),
		.mem_outb(mem_outb[22:27]));

	cb_mux_size48_mem mem_left_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_3_ccff_tail),
		.mem_out(mem_out[33:38]),
		.mem_outb(mem_outb[33:38]));

	cb_mux_size48_mem mem_left_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_4_ccff_tail),
		.mem_out(mem_out[44:49]),
		.mem_outb(mem_outb[44:49]));

	cb_mux_size48_mem mem_left_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_5_ccff_tail),
		.mem_out(mem_out[55:60]),
		.mem_outb(mem_outb[55:60]));

	cb_mux_size48_mem mem_left_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_6_ccff_tail),
		.mem_out(mem_out[66:71]),
		.mem_outb(mem_outb[66:71]));

	cb_mux_size48_mem mem_left_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_7_ccff_tail),
		.mem_out(mem_out[77:82]),
		.mem_outb(mem_outb[77:82]));

	cb_mux_size48_mem mem_left_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_8_ccff_tail),
		.mem_out(mem_out[94:99]),
		.mem_outb(mem_outb[94:99]));

	cb_mux_size48_mem mem_left_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_9_ccff_tail),
		.mem_out(mem_out[111:116]),
		.mem_outb(mem_outb[111:116]));

	cb_mux_size48_mem mem_left_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_10_ccff_tail),
		.mem_out(mem_out[128:133]),
		.mem_outb(mem_outb[128:133]));

	cb_mux_size48_mem mem_left_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_11_ccff_tail),
		.mem_out(mem_out[145:150]),
		.mem_outb(mem_outb[145:150]));

	cb_mux_size48_mem mem_left_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_12_ccff_tail),
		.mem_out(mem_out[162:167]),
		.mem_outb(mem_outb[162:167]));

	cb_mux_size48_mem mem_left_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_13_ccff_tail),
		.mem_out(mem_out[179:184]),
		.mem_outb(mem_outb[179:184]));

	cb_mux_size48_mem mem_left_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_14_ccff_tail),
		.mem_out(mem_out[196:201]),
		.mem_outb(mem_outb[196:201]));

	cb_mux_size48_mem mem_left_ipin_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_15_ccff_tail),
		.mem_out(mem_out[213:218]),
		.mem_outb(mem_outb[213:218]));

	cb_mux_size48_mem mem_right_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_29_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_16_ccff_tail),
		.mem_out(mem_out[434:439]),
		.mem_outb(mem_outb[434:439]));

	cb_mux_size48_mem mem_right_ipin_32 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_17_ccff_tail),
		.mem_out(mem_out[445:450]),
		.mem_outb(mem_outb[445:450]));

	cb_mux_size48_mem mem_right_ipin_35 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_18_ccff_tail),
		.mem_out(mem_out[462:467]),
		.mem_outb(mem_outb[462:467]));

	cb_mux_size48_mem mem_right_ipin_38 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size48_mem_19_ccff_tail),
		.mem_out(mem_out[479:484]),
		.mem_outb(mem_outb[479:484]));

	cb_mux_size16_mem mem_left_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_0_ccff_tail),
		.mem_out(mem_out[6:10]),
		.mem_outb(mem_outb[6:10]));

	cb_mux_size16_mem mem_left_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_1_ccff_tail),
		.mem_out(mem_out[17:21]),
		.mem_outb(mem_outb[17:21]));

	cb_mux_size16_mem mem_left_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_2_ccff_tail),
		.mem_out(mem_out[28:32]),
		.mem_outb(mem_outb[28:32]));

	cb_mux_size16_mem mem_left_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_3_ccff_tail),
		.mem_out(mem_out[39:43]),
		.mem_outb(mem_outb[39:43]));

	cb_mux_size16_mem mem_left_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_4_ccff_tail),
		.mem_out(mem_out[50:54]),
		.mem_outb(mem_outb[50:54]));

	cb_mux_size16_mem mem_left_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_5_ccff_tail),
		.mem_out(mem_out[61:65]),
		.mem_outb(mem_outb[61:65]));

	cb_mux_size16_mem mem_left_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_6_ccff_tail),
		.mem_out(mem_out[72:76]),
		.mem_outb(mem_outb[72:76]));

	cb_mux_size16_mem mem_left_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_7_ccff_tail),
		.mem_out(mem_out[83:87]),
		.mem_outb(mem_outb[83:87]));

	cb_mux_size16_mem mem_left_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_8_ccff_tail),
		.mem_out(mem_out[100:104]),
		.mem_outb(mem_outb[100:104]));

	cb_mux_size16_mem mem_left_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_9_ccff_tail),
		.mem_out(mem_out[117:121]),
		.mem_outb(mem_outb[117:121]));

	cb_mux_size16_mem mem_left_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_10_ccff_tail),
		.mem_out(mem_out[134:138]),
		.mem_outb(mem_outb[134:138]));

	cb_mux_size16_mem mem_left_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_11_ccff_tail),
		.mem_out(mem_out[151:155]),
		.mem_outb(mem_outb[151:155]));

	cb_mux_size16_mem mem_left_ipin_30 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_12_ccff_tail),
		.mem_out(mem_out[168:172]),
		.mem_outb(mem_outb[168:172]));

	cb_mux_size16_mem mem_left_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_13_ccff_tail),
		.mem_out(mem_out[185:189]),
		.mem_outb(mem_outb[185:189]));

	cb_mux_size16_mem mem_left_ipin_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_14_ccff_tail),
		.mem_out(mem_out[202:206]),
		.mem_outb(mem_outb[202:206]));

	cb_mux_size16_mem mem_left_ipin_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_15_ccff_tail),
		.mem_out(mem_out[219:223]),
		.mem_outb(mem_outb[219:223]));

	cb_mux_size16_mem mem_right_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_16_ccff_tail),
		.mem_out(mem_out[440:444]),
		.mem_outb(mem_outb[440:444]));

	cb_mux_size16_mem mem_right_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_17_ccff_tail),
		.mem_out(mem_out[457:461]),
		.mem_outb(mem_outb[457:461]));

	cb_mux_size16_mem mem_right_ipin_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_18_ccff_tail),
		.mem_out(mem_out[474:478]),
		.mem_outb(mem_outb[474:478]));

	cb_mux_size16_mem mem_right_ipin_40 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size56_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size16_mem_19_ccff_tail),
		.mem_out(mem_out[491:495]),
		.mem_outb(mem_outb[491:495]));

	cb_mux_size56_mem mem_left_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_0_ccff_tail),
		.mem_out(mem_out[88:93]),
		.mem_outb(mem_outb[88:93]));

	cb_mux_size56_mem mem_left_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_1_ccff_tail),
		.mem_out(mem_out[105:110]),
		.mem_outb(mem_outb[105:110]));

	cb_mux_size56_mem mem_left_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_2_ccff_tail),
		.mem_out(mem_out[122:127]),
		.mem_outb(mem_outb[122:127]));

	cb_mux_size56_mem mem_left_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_3_ccff_tail),
		.mem_out(mem_out[139:144]),
		.mem_outb(mem_outb[139:144]));

	cb_mux_size56_mem mem_left_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_4_ccff_tail),
		.mem_out(mem_out[156:161]),
		.mem_outb(mem_outb[156:161]));

	cb_mux_size56_mem mem_left_ipin_31 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_5_ccff_tail),
		.mem_out(mem_out[173:178]),
		.mem_outb(mem_outb[173:178]));

	cb_mux_size56_mem mem_left_ipin_34 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_6_ccff_tail),
		.mem_out(mem_out[190:195]),
		.mem_outb(mem_outb[190:195]));

	cb_mux_size56_mem mem_left_ipin_37 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_7_ccff_tail),
		.mem_out(mem_out[207:212]),
		.mem_outb(mem_outb[207:212]));

	cb_mux_size56_mem mem_right_ipin_33 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_8_ccff_tail),
		.mem_out(mem_out[451:456]),
		.mem_outb(mem_outb[451:456]));

	cb_mux_size56_mem mem_right_ipin_36 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_9_ccff_tail),
		.mem_out(mem_out[468:473]),
		.mem_outb(mem_outb[468:473]));

	cb_mux_size56_mem mem_right_ipin_39 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size48_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size56_mem_10_ccff_tail),
		.mem_out(mem_out[485:490]),
		.mem_outb(mem_outb[485:490]));

	cb_mux_size76_mem mem_right_ipin_0 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_0_ccff_tail),
		.mem_out(mem_out[224:230]),
		.mem_outb(mem_outb[224:230]));

	cb_mux_size76_mem mem_right_ipin_1 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_1_ccff_tail),
		.mem_out(mem_out[231:237]),
		.mem_outb(mem_outb[231:237]));

	cb_mux_size76_mem mem_right_ipin_2 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_2_ccff_tail),
		.mem_out(mem_out[238:244]),
		.mem_outb(mem_outb[238:244]));

	cb_mux_size76_mem mem_right_ipin_3 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_3_ccff_tail),
		.mem_out(mem_out[245:251]),
		.mem_outb(mem_outb[245:251]));

	cb_mux_size76_mem mem_right_ipin_4 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_4_ccff_tail),
		.mem_out(mem_out[252:258]),
		.mem_outb(mem_outb[252:258]));

	cb_mux_size76_mem mem_right_ipin_5 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_5_ccff_tail),
		.mem_out(mem_out[259:265]),
		.mem_outb(mem_outb[259:265]));

	cb_mux_size76_mem mem_right_ipin_6 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_6_ccff_tail),
		.mem_out(mem_out[266:272]),
		.mem_outb(mem_outb[266:272]));

	cb_mux_size76_mem mem_right_ipin_7 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_7_ccff_tail),
		.mem_out(mem_out[273:279]),
		.mem_outb(mem_outb[273:279]));

	cb_mux_size76_mem mem_right_ipin_8 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_8_ccff_tail),
		.mem_out(mem_out[280:286]),
		.mem_outb(mem_outb[280:286]));

	cb_mux_size76_mem mem_right_ipin_9 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_9_ccff_tail),
		.mem_out(mem_out[287:293]),
		.mem_outb(mem_outb[287:293]));

	cb_mux_size76_mem mem_right_ipin_10 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_10_ccff_tail),
		.mem_out(mem_out[294:300]),
		.mem_outb(mem_outb[294:300]));

	cb_mux_size76_mem mem_right_ipin_11 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_11_ccff_tail),
		.mem_out(mem_out[301:307]),
		.mem_outb(mem_outb[301:307]));

	cb_mux_size76_mem mem_right_ipin_12 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_12_ccff_tail),
		.mem_out(mem_out[308:314]),
		.mem_outb(mem_outb[308:314]));

	cb_mux_size76_mem mem_right_ipin_13 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_13_ccff_tail),
		.mem_out(mem_out[315:321]),
		.mem_outb(mem_outb[315:321]));

	cb_mux_size76_mem mem_right_ipin_14 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_14_ccff_tail),
		.mem_out(mem_out[322:328]),
		.mem_outb(mem_outb[322:328]));

	cb_mux_size76_mem mem_right_ipin_15 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_14_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_15_ccff_tail),
		.mem_out(mem_out[329:335]),
		.mem_outb(mem_outb[329:335]));

	cb_mux_size76_mem mem_right_ipin_16 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_15_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_16_ccff_tail),
		.mem_out(mem_out[336:342]),
		.mem_outb(mem_outb[336:342]));

	cb_mux_size76_mem mem_right_ipin_17 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_16_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_17_ccff_tail),
		.mem_out(mem_out[343:349]),
		.mem_outb(mem_outb[343:349]));

	cb_mux_size76_mem mem_right_ipin_18 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_17_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_18_ccff_tail),
		.mem_out(mem_out[350:356]),
		.mem_outb(mem_outb[350:356]));

	cb_mux_size76_mem mem_right_ipin_19 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_18_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_19_ccff_tail),
		.mem_out(mem_out[357:363]),
		.mem_outb(mem_outb[357:363]));

	cb_mux_size76_mem mem_right_ipin_20 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_20_ccff_tail),
		.mem_out(mem_out[364:370]),
		.mem_outb(mem_outb[364:370]));

	cb_mux_size76_mem mem_right_ipin_21 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_20_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_21_ccff_tail),
		.mem_out(mem_out[371:377]),
		.mem_outb(mem_outb[371:377]));

	cb_mux_size76_mem mem_right_ipin_22 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_21_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_22_ccff_tail),
		.mem_out(mem_out[378:384]),
		.mem_outb(mem_outb[378:384]));

	cb_mux_size76_mem mem_right_ipin_23 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_22_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_23_ccff_tail),
		.mem_out(mem_out[385:391]),
		.mem_outb(mem_outb[385:391]));

	cb_mux_size76_mem mem_right_ipin_24 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_23_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_24_ccff_tail),
		.mem_out(mem_out[392:398]),
		.mem_outb(mem_outb[392:398]));

	cb_mux_size76_mem mem_right_ipin_25 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_24_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_25_ccff_tail),
		.mem_out(mem_out[399:405]),
		.mem_outb(mem_outb[399:405]));

	cb_mux_size76_mem mem_right_ipin_26 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_25_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_26_ccff_tail),
		.mem_out(mem_out[406:412]),
		.mem_outb(mem_outb[406:412]));

	cb_mux_size76_mem mem_right_ipin_27 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_26_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_27_ccff_tail),
		.mem_out(mem_out[413:419]),
		.mem_outb(mem_outb[413:419]));

	cb_mux_size76_mem mem_right_ipin_28 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_27_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_28_ccff_tail),
		.mem_out(mem_out[420:426]),
		.mem_outb(mem_outb[420:426]));

	cb_mux_size76_mem mem_right_ipin_29 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size76_mem_28_ccff_tail),
		.ccff_tail(cb_mux_size76_mem_29_ccff_tail),
		.mem_out(mem_out[427:433]),
		.mem_outb(mem_outb[427:433]));

	cb_mux_size8_mem mem_right_ipin_41 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size16_mem_19_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_0_ccff_tail),
		.mem_out(mem_out[496:499]),
		.mem_outb(mem_outb[496:499]));

	cb_mux_size8_mem mem_right_ipin_42 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_0_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_1_ccff_tail),
		.mem_out(mem_out[500:503]),
		.mem_outb(mem_outb[500:503]));

	cb_mux_size8_mem mem_right_ipin_43 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_1_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_2_ccff_tail),
		.mem_out(mem_out[504:507]),
		.mem_outb(mem_outb[504:507]));

	cb_mux_size8_mem mem_right_ipin_44 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_2_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_3_ccff_tail),
		.mem_out(mem_out[508:511]),
		.mem_outb(mem_outb[508:511]));

	cb_mux_size8_mem mem_right_ipin_45 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_3_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_4_ccff_tail),
		.mem_out(mem_out[512:515]),
		.mem_outb(mem_outb[512:515]));

	cb_mux_size8_mem mem_right_ipin_46 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_4_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_5_ccff_tail),
		.mem_out(mem_out[516:519]),
		.mem_outb(mem_outb[516:519]));

	cb_mux_size8_mem mem_right_ipin_47 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_5_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_6_ccff_tail),
		.mem_out(mem_out[520:523]),
		.mem_outb(mem_outb[520:523]));

	cb_mux_size8_mem mem_right_ipin_48 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_6_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_7_ccff_tail),
		.mem_out(mem_out[524:527]),
		.mem_outb(mem_outb[524:527]));

	cb_mux_size8_mem mem_right_ipin_49 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_7_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_8_ccff_tail),
		.mem_out(mem_out[528:531]),
		.mem_outb(mem_outb[528:531]));

	cb_mux_size8_mem mem_right_ipin_50 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_8_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_9_ccff_tail),
		.mem_out(mem_out[532:535]),
		.mem_outb(mem_outb[532:535]));

	cb_mux_size8_mem mem_right_ipin_51 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_9_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_10_ccff_tail),
		.mem_out(mem_out[536:539]),
		.mem_outb(mem_outb[536:539]));

	cb_mux_size8_mem mem_right_ipin_52 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_10_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_11_ccff_tail),
		.mem_out(mem_out[540:543]),
		.mem_outb(mem_outb[540:543]));

	cb_mux_size8_mem mem_right_ipin_53 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_11_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_12_ccff_tail),
		.mem_out(mem_out[544:547]),
		.mem_outb(mem_outb[544:547]));

	cb_mux_size8_mem mem_right_ipin_54 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_12_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_13_ccff_tail),
		.mem_out(mem_out[548:551]),
		.mem_outb(mem_outb[548:551]));

	cb_mux_size8_mem mem_right_ipin_55 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_13_ccff_tail),
		.ccff_tail(cb_mux_size8_mem_14_ccff_tail),
		.mem_out(mem_out[552:555]),
		.mem_outb(mem_outb[552:555]));

	cb_mux_size8_mem mem_right_ipin_56 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(cb_mux_size8_mem_14_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mem_out[556:559]),
		.mem_outb(mem_outb[556:559]));

endmodule
// ----- END Verilog module for cby_6__config_group_mem_size560 -----




