//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//-------------------------------------------
// ----- Verilog module for sb_0_ -----
module sb_0_(config_enable,
             prog_reset,
             prog_clk,
             chany_top_in,
             top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_,
             top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_,
             chanx_right_in,
             right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_,
             right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_,
             chany_bottom_in,
             chanx_left_in,
             ccff_head,
             chany_top_out,
             chanx_right_out,
             chany_bottom_out,
             chanx_left_out,
             ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] config_enable;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:63] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:63] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_;
//----- INPUT PORTS -----
input [0:31] chany_bottom_in;
//----- INPUT PORTS -----
input [0:63] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:63] chany_top_out;
//----- OUTPUT PORTS -----
output [0:63] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:31] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:63] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] clk_mux_size3_0_sram;
wire [0:1] clk_mux_size3_0_sram_inv;
wire [0:1] clk_mux_size3_10_sram;
wire [0:1] clk_mux_size3_10_sram_inv;
wire [0:1] clk_mux_size3_11_sram;
wire [0:1] clk_mux_size3_11_sram_inv;
wire [0:1] clk_mux_size3_12_sram;
wire [0:1] clk_mux_size3_12_sram_inv;
wire [0:1] clk_mux_size3_13_sram;
wire [0:1] clk_mux_size3_13_sram_inv;
wire [0:1] clk_mux_size3_14_sram;
wire [0:1] clk_mux_size3_14_sram_inv;
wire [0:1] clk_mux_size3_15_sram;
wire [0:1] clk_mux_size3_15_sram_inv;
wire [0:1] clk_mux_size3_16_sram;
wire [0:1] clk_mux_size3_16_sram_inv;
wire [0:1] clk_mux_size3_17_sram;
wire [0:1] clk_mux_size3_17_sram_inv;
wire [0:1] clk_mux_size3_18_sram;
wire [0:1] clk_mux_size3_18_sram_inv;
wire [0:1] clk_mux_size3_19_sram;
wire [0:1] clk_mux_size3_19_sram_inv;
wire [0:1] clk_mux_size3_1_sram;
wire [0:1] clk_mux_size3_1_sram_inv;
wire [0:1] clk_mux_size3_20_sram;
wire [0:1] clk_mux_size3_20_sram_inv;
wire [0:1] clk_mux_size3_21_sram;
wire [0:1] clk_mux_size3_21_sram_inv;
wire [0:1] clk_mux_size3_22_sram;
wire [0:1] clk_mux_size3_22_sram_inv;
wire [0:1] clk_mux_size3_23_sram;
wire [0:1] clk_mux_size3_23_sram_inv;
wire [0:1] clk_mux_size3_24_sram;
wire [0:1] clk_mux_size3_24_sram_inv;
wire [0:1] clk_mux_size3_25_sram;
wire [0:1] clk_mux_size3_25_sram_inv;
wire [0:1] clk_mux_size3_26_sram;
wire [0:1] clk_mux_size3_26_sram_inv;
wire [0:1] clk_mux_size3_27_sram;
wire [0:1] clk_mux_size3_27_sram_inv;
wire [0:1] clk_mux_size3_28_sram;
wire [0:1] clk_mux_size3_28_sram_inv;
wire [0:1] clk_mux_size3_29_sram;
wire [0:1] clk_mux_size3_29_sram_inv;
wire [0:1] clk_mux_size3_2_sram;
wire [0:1] clk_mux_size3_2_sram_inv;
wire [0:1] clk_mux_size3_30_sram;
wire [0:1] clk_mux_size3_30_sram_inv;
wire [0:1] clk_mux_size3_31_sram;
wire [0:1] clk_mux_size3_31_sram_inv;
wire [0:1] clk_mux_size3_32_sram;
wire [0:1] clk_mux_size3_32_sram_inv;
wire [0:1] clk_mux_size3_33_sram;
wire [0:1] clk_mux_size3_33_sram_inv;
wire [0:1] clk_mux_size3_34_sram;
wire [0:1] clk_mux_size3_34_sram_inv;
wire [0:1] clk_mux_size3_35_sram;
wire [0:1] clk_mux_size3_35_sram_inv;
wire [0:1] clk_mux_size3_36_sram;
wire [0:1] clk_mux_size3_36_sram_inv;
wire [0:1] clk_mux_size3_37_sram;
wire [0:1] clk_mux_size3_37_sram_inv;
wire [0:1] clk_mux_size3_38_sram;
wire [0:1] clk_mux_size3_38_sram_inv;
wire [0:1] clk_mux_size3_39_sram;
wire [0:1] clk_mux_size3_39_sram_inv;
wire [0:1] clk_mux_size3_3_sram;
wire [0:1] clk_mux_size3_3_sram_inv;
wire [0:1] clk_mux_size3_40_sram;
wire [0:1] clk_mux_size3_40_sram_inv;
wire [0:1] clk_mux_size3_41_sram;
wire [0:1] clk_mux_size3_41_sram_inv;
wire [0:1] clk_mux_size3_42_sram;
wire [0:1] clk_mux_size3_42_sram_inv;
wire [0:1] clk_mux_size3_43_sram;
wire [0:1] clk_mux_size3_43_sram_inv;
wire [0:1] clk_mux_size3_44_sram;
wire [0:1] clk_mux_size3_44_sram_inv;
wire [0:1] clk_mux_size3_45_sram;
wire [0:1] clk_mux_size3_45_sram_inv;
wire [0:1] clk_mux_size3_46_sram;
wire [0:1] clk_mux_size3_46_sram_inv;
wire [0:1] clk_mux_size3_47_sram;
wire [0:1] clk_mux_size3_47_sram_inv;
wire [0:1] clk_mux_size3_48_sram;
wire [0:1] clk_mux_size3_48_sram_inv;
wire [0:1] clk_mux_size3_49_sram;
wire [0:1] clk_mux_size3_49_sram_inv;
wire [0:1] clk_mux_size3_4_sram;
wire [0:1] clk_mux_size3_4_sram_inv;
wire [0:1] clk_mux_size3_50_sram;
wire [0:1] clk_mux_size3_50_sram_inv;
wire [0:1] clk_mux_size3_51_sram;
wire [0:1] clk_mux_size3_51_sram_inv;
wire [0:1] clk_mux_size3_52_sram;
wire [0:1] clk_mux_size3_52_sram_inv;
wire [0:1] clk_mux_size3_53_sram;
wire [0:1] clk_mux_size3_53_sram_inv;
wire [0:1] clk_mux_size3_54_sram;
wire [0:1] clk_mux_size3_54_sram_inv;
wire [0:1] clk_mux_size3_55_sram;
wire [0:1] clk_mux_size3_55_sram_inv;
wire [0:1] clk_mux_size3_56_sram;
wire [0:1] clk_mux_size3_56_sram_inv;
wire [0:1] clk_mux_size3_57_sram;
wire [0:1] clk_mux_size3_57_sram_inv;
wire [0:1] clk_mux_size3_58_sram;
wire [0:1] clk_mux_size3_58_sram_inv;
wire [0:1] clk_mux_size3_59_sram;
wire [0:1] clk_mux_size3_59_sram_inv;
wire [0:1] clk_mux_size3_5_sram;
wire [0:1] clk_mux_size3_5_sram_inv;
wire [0:1] clk_mux_size3_60_sram;
wire [0:1] clk_mux_size3_60_sram_inv;
wire [0:1] clk_mux_size3_61_sram;
wire [0:1] clk_mux_size3_61_sram_inv;
wire [0:1] clk_mux_size3_62_sram;
wire [0:1] clk_mux_size3_62_sram_inv;
wire [0:1] clk_mux_size3_63_sram;
wire [0:1] clk_mux_size3_63_sram_inv;
wire [0:1] clk_mux_size3_6_sram;
wire [0:1] clk_mux_size3_6_sram_inv;
wire [0:1] clk_mux_size3_7_sram;
wire [0:1] clk_mux_size3_7_sram_inv;
wire [0:1] clk_mux_size3_8_sram;
wire [0:1] clk_mux_size3_8_sram_inv;
wire [0:1] clk_mux_size3_9_sram;
wire [0:1] clk_mux_size3_9_sram_inv;
wire [0:264] sb_0__config_group_mem_size265_0_mem_out;
wire [0:264] sb_0__config_group_mem_size265_0_mem_outb;
wire [0:1] sb_mux_size2_0_sram;
wire [0:1] sb_mux_size2_0_sram_inv;
wire [0:1] sb_mux_size2_1_sram;
wire [0:1] sb_mux_size2_1_sram_inv;
wire [0:1] sb_mux_size3_0_sram;
wire [0:1] sb_mux_size3_0_sram_inv;
wire [0:1] sb_mux_size3_1_sram;
wire [0:1] sb_mux_size3_1_sram_inv;
wire [0:1] sb_mux_size3_2_sram;
wire [0:1] sb_mux_size3_2_sram_inv;
wire [0:1] sb_mux_size3_3_sram;
wire [0:1] sb_mux_size3_3_sram_inv;
wire [0:1] sb_mux_size3_4_sram;
wire [0:1] sb_mux_size3_4_sram_inv;
wire [0:2] sb_mux_size4_0_sram;
wire [0:2] sb_mux_size4_0_sram_inv;
wire [0:2] sb_mux_size4_10_sram;
wire [0:2] sb_mux_size4_10_sram_inv;
wire [0:2] sb_mux_size4_11_sram;
wire [0:2] sb_mux_size4_11_sram_inv;
wire [0:2] sb_mux_size4_12_sram;
wire [0:2] sb_mux_size4_12_sram_inv;
wire [0:2] sb_mux_size4_13_sram;
wire [0:2] sb_mux_size4_13_sram_inv;
wire [0:2] sb_mux_size4_14_sram;
wire [0:2] sb_mux_size4_14_sram_inv;
wire [0:2] sb_mux_size4_15_sram;
wire [0:2] sb_mux_size4_15_sram_inv;
wire [0:2] sb_mux_size4_1_sram;
wire [0:2] sb_mux_size4_1_sram_inv;
wire [0:2] sb_mux_size4_2_sram;
wire [0:2] sb_mux_size4_2_sram_inv;
wire [0:2] sb_mux_size4_3_sram;
wire [0:2] sb_mux_size4_3_sram_inv;
wire [0:2] sb_mux_size4_4_sram;
wire [0:2] sb_mux_size4_4_sram_inv;
wire [0:2] sb_mux_size4_5_sram;
wire [0:2] sb_mux_size4_5_sram_inv;
wire [0:2] sb_mux_size4_6_sram;
wire [0:2] sb_mux_size4_6_sram_inv;
wire [0:2] sb_mux_size4_7_sram;
wire [0:2] sb_mux_size4_7_sram_inv;
wire [0:2] sb_mux_size4_8_sram;
wire [0:2] sb_mux_size4_8_sram_inv;
wire [0:2] sb_mux_size4_9_sram;
wire [0:2] sb_mux_size4_9_sram_inv;
wire [0:2] sb_mux_size5_0_sram;
wire [0:2] sb_mux_size5_0_sram_inv;
wire [0:2] sb_mux_size5_10_sram;
wire [0:2] sb_mux_size5_10_sram_inv;
wire [0:2] sb_mux_size5_11_sram;
wire [0:2] sb_mux_size5_11_sram_inv;
wire [0:2] sb_mux_size5_12_sram;
wire [0:2] sb_mux_size5_12_sram_inv;
wire [0:2] sb_mux_size5_13_sram;
wire [0:2] sb_mux_size5_13_sram_inv;
wire [0:2] sb_mux_size5_14_sram;
wire [0:2] sb_mux_size5_14_sram_inv;
wire [0:2] sb_mux_size5_15_sram;
wire [0:2] sb_mux_size5_15_sram_inv;
wire [0:2] sb_mux_size5_16_sram;
wire [0:2] sb_mux_size5_16_sram_inv;
wire [0:2] sb_mux_size5_1_sram;
wire [0:2] sb_mux_size5_1_sram_inv;
wire [0:2] sb_mux_size5_2_sram;
wire [0:2] sb_mux_size5_2_sram_inv;
wire [0:2] sb_mux_size5_3_sram;
wire [0:2] sb_mux_size5_3_sram_inv;
wire [0:2] sb_mux_size5_4_sram;
wire [0:2] sb_mux_size5_4_sram_inv;
wire [0:2] sb_mux_size5_5_sram;
wire [0:2] sb_mux_size5_5_sram_inv;
wire [0:2] sb_mux_size5_6_sram;
wire [0:2] sb_mux_size5_6_sram_inv;
wire [0:2] sb_mux_size5_7_sram;
wire [0:2] sb_mux_size5_7_sram_inv;
wire [0:2] sb_mux_size5_8_sram;
wire [0:2] sb_mux_size5_8_sram_inv;
wire [0:2] sb_mux_size5_9_sram;
wire [0:2] sb_mux_size5_9_sram_inv;
wire [0:2] sb_mux_size6_0_sram;
wire [0:2] sb_mux_size6_0_sram_inv;
wire [0:2] sb_mux_size6_1_sram;
wire [0:2] sb_mux_size6_1_sram_inv;
wire [0:2] sb_mux_size6_2_sram;
wire [0:2] sb_mux_size6_2_sram_inv;
wire [0:2] sb_mux_size6_3_sram;
wire [0:2] sb_mux_size6_3_sram_inv;
wire [0:2] sb_mux_size6_4_sram;
wire [0:2] sb_mux_size6_4_sram_inv;
wire [0:2] sb_mux_size6_5_sram;
wire [0:2] sb_mux_size6_5_sram_inv;
wire [0:2] sb_mux_size6_6_sram;
wire [0:2] sb_mux_size6_6_sram_inv;
wire [0:2] sb_mux_size6_7_sram;
wire [0:2] sb_mux_size6_7_sram_inv;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chany_top_out[18] = top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_[0];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[32] = chanx_right_in[32];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[33];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[34];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[35];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[36] = chanx_right_in[36];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[37];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[38];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[39];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[40] = chanx_right_in[40];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[41];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[42];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[43];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[44] = chanx_right_in[44];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[45];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[46];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[47];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[48] = chanx_right_in[48];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[49];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[50];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[51];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[52] = chanx_right_in[52];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[53];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[54];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[55];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[56] = chanx_right_in[56];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[57];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[58];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[59];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[60] = chanx_right_in[60];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[61];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[62];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[63];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chanx_left_in[2];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chanx_left_in[3];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[28] = chanx_left_in[4];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chanx_left_in[5];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chanx_left_in[7];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chanx_left_in[9];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[24] = chanx_left_in[11];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chanx_left_in[15];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chanx_left_in[19];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chanx_left_in[23];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[20] = chanx_left_in[27];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[32] = chanx_left_in[32];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[33];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[34];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[35];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[36] = chanx_left_in[36];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[37];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[38];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[39];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[40] = chanx_left_in[40];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[41];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[42];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[43];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[44] = chanx_left_in[44];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[45];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[46];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[47];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[48] = chanx_left_in[48];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[49];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[50];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[51];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[52] = chanx_left_in[52];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[53];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[54];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[55];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[56] = chanx_left_in[56];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[57];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[58];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[59];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[60] = chanx_left_in[60];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[61];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[62];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[63];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	sb_mux_size6 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[1], chanx_right_in[6], chanx_left_in[0], chanx_left_in[6]}),
		.sram(sb_mux_size6_0_sram[0:2]),
		.sram_inv(sb_mux_size6_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	sb_mux_size6 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[14], chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[1]}),
		.sram(sb_mux_size6_1_sram[0:2]),
		.sram_inv(sb_mux_size6_1_sram_inv[0:2]),
		.out(chanx_right_out[1]));

	sb_mux_size6 mux_right_track_12 (
		.in({chany_top_in[5], chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[7]}),
		.sram(sb_mux_size6_2_sram[0:2]),
		.sram_inv(sb_mux_size6_2_sram_inv[0:2]),
		.out(chanx_right_out[6]));

	sb_mux_size6 mux_right_track_16 (
		.in({chany_top_in[6], chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[9]}),
		.sram(sb_mux_size6_3_sram[0:2]),
		.sram_inv(sb_mux_size6_3_sram_inv[0:2]),
		.out(chanx_right_out[8]));

	sb_mux_size6 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[14], chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[0]}),
		.sram(sb_mux_size6_4_sram[0:2]),
		.sram_inv(sb_mux_size6_4_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	sb_mux_size6 mux_left_track_13 (
		.in({chany_top_in[8], chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[7]}),
		.sram(sb_mux_size6_5_sram[0:2]),
		.sram_inv(sb_mux_size6_5_sram_inv[0:2]),
		.out(chanx_left_out[6]));

	sb_mux_size6 mux_left_track_17 (
		.in({chany_top_in[7], chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[9]}),
		.sram(sb_mux_size6_6_sram[0:2]),
		.sram_inv(sb_mux_size6_6_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	sb_mux_size6 mux_left_track_41 (
		.in({chany_top_in[3], chany_top_in[17], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[23]}),
		.sram(sb_mux_size6_7_sram[0:2]),
		.sram_inv(sb_mux_size6_7_sram_inv[0:2]),
		.out(chanx_left_out[20]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_top_track_0 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[0:2]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[0:2]),
		.mem_out(sb_mux_size6_0_sram[0:2]),
		.mem_outb(sb_mux_size6_0_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_right_track_2 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[120:122]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[120:122]),
		.mem_out(sb_mux_size6_1_sram[0:2]),
		.mem_outb(sb_mux_size6_1_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_right_track_12 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[135:137]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[135:137]),
		.mem_out(sb_mux_size6_2_sram[0:2]),
		.mem_outb(sb_mux_size6_2_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_right_track_16 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[138:140]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[138:140]),
		.mem_out(sb_mux_size6_3_sram[0:2]),
		.mem_outb(sb_mux_size6_3_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_left_track_1 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[223:225]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[223:225]),
		.mem_out(sb_mux_size6_4_sram[0:2]),
		.mem_outb(sb_mux_size6_4_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_left_track_13 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[241:243]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[241:243]),
		.mem_out(sb_mux_size6_5_sram[0:2]),
		.mem_outb(sb_mux_size6_5_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_left_track_17 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[244:246]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[244:246]),
		.mem_out(sb_mux_size6_6_sram[0:2]),
		.mem_outb(sb_mux_size6_6_sram_inv[0:2]));

	sb_mux_size6_feedthrough_mem feedthrough_mem_left_track_41 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[256:258]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[256:258]),
		.mem_out(sb_mux_size6_7_sram[0:2]),
		.mem_outb(sb_mux_size6_7_sram_inv[0:2]));

	sb_mux_size5 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[2], chanx_right_in[8], chanx_left_in[8]}),
		.sram(sb_mux_size5_0_sram[0:2]),
		.sram_inv(sb_mux_size5_0_sram_inv[0:2]),
		.out(chany_top_out[1]));

	sb_mux_size5 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[9], chanx_right_in[16], chanx_left_in[16]}),
		.sram(sb_mux_size5_1_sram[0:2]),
		.sram_inv(sb_mux_size5_1_sram_inv[0:2]),
		.out(chany_top_out[6]));

	sb_mux_size5 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[11], chanx_right_in[17], chanx_left_in[17]}),
		.sram(sb_mux_size5_2_sram[0:2]),
		.sram_inv(sb_mux_size5_2_sram_inv[0:2]),
		.out(chany_top_out[7]));

	sb_mux_size5 mux_right_track_0 (
		.in({chany_top_in[13], chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[0]}),
		.sram(sb_mux_size5_3_sram[0:2]),
		.sram_inv(sb_mux_size5_3_sram_inv[0:2]),
		.out(chanx_right_out[0]));

	sb_mux_size5 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[15], chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_left_in[2]}),
		.sram(sb_mux_size5_4_sram[0:2]),
		.sram_inv(sb_mux_size5_4_sram_inv[0:2]),
		.out(chanx_right_out[2]));

	sb_mux_size5 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[16], chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_left_in[3]}),
		.sram(sb_mux_size5_5_sram[0:2]),
		.sram_inv(sb_mux_size5_5_sram_inv[0:2]),
		.out(chanx_right_out[3]));

	sb_mux_size5 mux_right_track_8 (
		.in({chany_top_in[3], chany_top_in[17], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_left_in[4]}),
		.sram(sb_mux_size5_6_sram[0:2]),
		.sram_inv(sb_mux_size5_6_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	sb_mux_size5 mux_right_track_20 (
		.in({chany_top_in[7], chany_top_in[21], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[11]}),
		.sram(sb_mux_size5_7_sram[0:2]),
		.sram_inv(sb_mux_size5_7_sram_inv[0:2]),
		.out(chanx_right_out[10]));

	sb_mux_size5 mux_right_track_24 (
		.in({chany_top_in[8], chany_top_in[22], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[15]}),
		.sram(sb_mux_size5_8_sram[0:2]),
		.sram_inv(sb_mux_size5_8_sram_inv[0:2]),
		.out(chanx_right_out[12]));

	sb_mux_size5 mux_right_track_32 (
		.in({chany_top_in[9], chany_top_in[23], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_left_in[19]}),
		.sram(sb_mux_size5_9_sram[0:2]),
		.sram_inv(sb_mux_size5_9_sram_inv[0:2]),
		.out(chanx_right_out[16]));

	sb_mux_size5 mux_right_track_40 (
		.in({chany_top_in[10], chany_top_in[24], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[23]}),
		.sram(sb_mux_size5_10_sram[0:2]),
		.sram_inv(sb_mux_size5_10_sram_inv[0:2]),
		.out(chanx_right_out[20]));

	sb_mux_size5 mux_left_track_3 (
		.in({chany_top_in[13], chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_right_in[1]}),
		.sram(sb_mux_size5_11_sram[0:2]),
		.sram_inv(sb_mux_size5_11_sram_inv[0:2]),
		.out(chanx_left_out[1]));

	sb_mux_size5 mux_left_track_21 (
		.in({chany_top_in[6], chany_top_in[20], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[11]}),
		.sram(sb_mux_size5_12_sram[0:2]),
		.sram_inv(sb_mux_size5_12_sram_inv[0:2]),
		.out(chanx_left_out[10]));

	sb_mux_size5 mux_left_track_25 (
		.in({chany_top_in[5], chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_0__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[15]}),
		.sram(sb_mux_size5_13_sram[0:2]),
		.sram_inv(sb_mux_size5_13_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	sb_mux_size5 mux_left_track_33 (
		.in({chany_top_in[4], chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_1__pin_a2f_o_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_a2f_o_0_, chanx_right_in[19]}),
		.sram(sb_mux_size5_14_sram[0:2]),
		.sram_inv(sb_mux_size5_14_sram_inv[0:2]),
		.out(chanx_left_out[16]));

	sb_mux_size5 mux_left_track_49 (
		.in({chany_top_in[2], chany_top_in[16], chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[27]}),
		.sram(sb_mux_size5_15_sram[0:2]),
		.sram_inv(sb_mux_size5_15_sram_inv[0:2]),
		.out(chanx_left_out[24]));

	sb_mux_size5 mux_left_track_57 (
		.in({chany_top_in[1], chany_top_in[15], chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[31]}),
		.sram(sb_mux_size5_16_sram[0:2]),
		.sram_inv(sb_mux_size5_16_sram_inv[0:2]),
		.out(chanx_left_out[28]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_top_track_2 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[3:5]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[3:5]),
		.mem_out(sb_mux_size5_0_sram[0:2]),
		.mem_outb(sb_mux_size5_0_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_top_track_12 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[18:20]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[18:20]),
		.mem_out(sb_mux_size5_1_sram[0:2]),
		.mem_outb(sb_mux_size5_1_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_top_track_14 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[21:23]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[21:23]),
		.mem_out(sb_mux_size5_2_sram[0:2]),
		.mem_outb(sb_mux_size5_2_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_0 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[117:119]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[117:119]),
		.mem_out(sb_mux_size5_3_sram[0:2]),
		.mem_outb(sb_mux_size5_3_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_4 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[123:125]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[123:125]),
		.mem_out(sb_mux_size5_4_sram[0:2]),
		.mem_outb(sb_mux_size5_4_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_6 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[126:128]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[126:128]),
		.mem_out(sb_mux_size5_5_sram[0:2]),
		.mem_outb(sb_mux_size5_5_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_8 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[129:131]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[129:131]),
		.mem_out(sb_mux_size5_6_sram[0:2]),
		.mem_outb(sb_mux_size5_6_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_20 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[141:143]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[141:143]),
		.mem_out(sb_mux_size5_7_sram[0:2]),
		.mem_outb(sb_mux_size5_7_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_24 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[144:146]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[144:146]),
		.mem_out(sb_mux_size5_8_sram[0:2]),
		.mem_outb(sb_mux_size5_8_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_32 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[147:149]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[147:149]),
		.mem_out(sb_mux_size5_9_sram[0:2]),
		.mem_outb(sb_mux_size5_9_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_right_track_40 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[150:152]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[150:152]),
		.mem_out(sb_mux_size5_10_sram[0:2]),
		.mem_outb(sb_mux_size5_10_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_3 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[226:228]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[226:228]),
		.mem_out(sb_mux_size5_11_sram[0:2]),
		.mem_outb(sb_mux_size5_11_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_21 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[247:249]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[247:249]),
		.mem_out(sb_mux_size5_12_sram[0:2]),
		.mem_outb(sb_mux_size5_12_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_25 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[250:252]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[250:252]),
		.mem_out(sb_mux_size5_13_sram[0:2]),
		.mem_outb(sb_mux_size5_13_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_33 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[253:255]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[253:255]),
		.mem_out(sb_mux_size5_14_sram[0:2]),
		.mem_outb(sb_mux_size5_14_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_49 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[259:261]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[259:261]),
		.mem_out(sb_mux_size5_15_sram[0:2]),
		.mem_outb(sb_mux_size5_15_sram_inv[0:2]));

	sb_mux_size5_feedthrough_mem feedthrough_mem_left_track_57 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[262:264]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[262:264]),
		.mem_out(sb_mux_size5_16_sram[0:2]),
		.mem_outb(sb_mux_size5_16_sram_inv[0:2]));

	sb_mux_size4 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_right_in[3], chanx_right_in[10], chanx_left_in[10]}),
		.sram(sb_mux_size4_0_sram[0:2]),
		.sram_inv(sb_mux_size4_0_sram_inv[0:2]),
		.out(chany_top_out[2]));

	sb_mux_size4 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[4], chanx_right_in[12], chanx_left_in[12]}),
		.sram(sb_mux_size4_1_sram[0:2]),
		.sram_inv(sb_mux_size4_1_sram_inv[0:2]),
		.out(chany_top_out[3]));

	sb_mux_size4 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[5], chanx_right_in[13], chanx_left_in[13]}),
		.sram(sb_mux_size4_2_sram[0:2]),
		.sram_inv(sb_mux_size4_2_sram_inv[0:2]),
		.out(chany_top_out[4]));

	sb_mux_size4 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[7], chanx_right_in[14], chanx_left_in[14]}),
		.sram(sb_mux_size4_3_sram[0:2]),
		.sram_inv(sb_mux_size4_3_sram_inv[0:2]),
		.out(chany_top_out[5]));

	sb_mux_size4 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_right_in[15], chanx_right_in[18], chanx_left_in[18]}),
		.sram(sb_mux_size4_4_sram[0:2]),
		.sram_inv(sb_mux_size4_4_sram_inv[0:2]),
		.out(chany_top_out[8]));

	sb_mux_size4 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[19:20], chanx_left_in[20]}),
		.sram(sb_mux_size4_5_sram[0:2]),
		.sram_inv(sb_mux_size4_5_sram_inv[0:2]),
		.out(chany_top_out[9]));

	sb_mux_size4 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[21], chanx_right_in[23], chanx_left_in[21]}),
		.sram(sb_mux_size4_6_sram[0:2]),
		.sram_inv(sb_mux_size4_6_sram_inv[0:2]),
		.out(chany_top_out[10]));

	sb_mux_size4 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[22], chanx_right_in[27], chanx_left_in[22]}),
		.sram(sb_mux_size4_7_sram[0:2]),
		.sram_inv(sb_mux_size4_7_sram_inv[0:2]),
		.out(chany_top_out[11]));

	sb_mux_size4 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_a2f_o_0_, chanx_right_in[24], chanx_right_in[31], chanx_left_in[24]}),
		.sram(sb_mux_size4_8_sram[0:2]),
		.sram_inv(sb_mux_size4_8_sram_inv[0:2]),
		.out(chany_top_out[12]));

	sb_mux_size4 mux_right_track_10 (
		.in({chany_top_in[4], chany_top_in[18], right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_left_in[5]}),
		.sram(sb_mux_size4_9_sram[0:2]),
		.sram_inv(sb_mux_size4_9_sram_inv[0:2]),
		.out(chanx_right_out[5]));

	sb_mux_size4 mux_right_track_48 (
		.in({chany_top_in[11], chany_top_in[25], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_left_in[27]}),
		.sram(sb_mux_size4_10_sram[0:2]),
		.sram_inv(sb_mux_size4_10_sram_inv[0:2]),
		.out(chanx_right_out[24]));

	sb_mux_size4 mux_right_track_56 (
		.in({chany_top_in[12], chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_left_in[31]}),
		.sram(sb_mux_size4_11_sram[0:2]),
		.sram_inv(sb_mux_size4_11_sram_inv[0:2]),
		.out(chanx_right_out[28]));

	sb_mux_size4 mux_left_track_5 (
		.in({chany_top_in[12], chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_right_in[2]}),
		.sram(sb_mux_size4_12_sram[0:2]),
		.sram_inv(sb_mux_size4_12_sram_inv[0:2]),
		.out(chanx_left_out[2]));

	sb_mux_size4 mux_left_track_7 (
		.in({chany_top_in[11], chany_top_in[25], right_bottom_grid_top_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[3]}),
		.sram(sb_mux_size4_13_sram[0:2]),
		.sram_inv(sb_mux_size4_13_sram_inv[0:2]),
		.out(chanx_left_out[3]));

	sb_mux_size4 mux_left_track_9 (
		.in({chany_top_in[10], chany_top_in[24], right_bottom_grid_top_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[4]}),
		.sram(sb_mux_size4_14_sram[0:2]),
		.sram_inv(sb_mux_size4_14_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	sb_mux_size4 mux_left_track_11 (
		.in({chany_top_in[9], chany_top_in[23], right_bottom_grid_top_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[5]}),
		.sram(sb_mux_size4_15_sram[0:2]),
		.sram_inv(sb_mux_size4_15_sram_inv[0:2]),
		.out(chanx_left_out[5]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_4 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[6:8]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[6:8]),
		.mem_out(sb_mux_size4_0_sram[0:2]),
		.mem_outb(sb_mux_size4_0_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_6 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[9:11]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[9:11]),
		.mem_out(sb_mux_size4_1_sram[0:2]),
		.mem_outb(sb_mux_size4_1_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_8 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[12:14]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[12:14]),
		.mem_out(sb_mux_size4_2_sram[0:2]),
		.mem_outb(sb_mux_size4_2_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_10 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[15:17]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[15:17]),
		.mem_out(sb_mux_size4_3_sram[0:2]),
		.mem_outb(sb_mux_size4_3_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_16 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[24:26]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[24:26]),
		.mem_out(sb_mux_size4_4_sram[0:2]),
		.mem_outb(sb_mux_size4_4_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_18 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[27:29]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[27:29]),
		.mem_out(sb_mux_size4_5_sram[0:2]),
		.mem_outb(sb_mux_size4_5_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_20 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[30:32]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[30:32]),
		.mem_out(sb_mux_size4_6_sram[0:2]),
		.mem_outb(sb_mux_size4_6_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_22 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[33:35]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[33:35]),
		.mem_out(sb_mux_size4_7_sram[0:2]),
		.mem_outb(sb_mux_size4_7_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_top_track_24 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[36:38]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[36:38]),
		.mem_out(sb_mux_size4_8_sram[0:2]),
		.mem_outb(sb_mux_size4_8_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_right_track_10 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[132:134]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[132:134]),
		.mem_out(sb_mux_size4_9_sram[0:2]),
		.mem_outb(sb_mux_size4_9_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_right_track_48 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[153:155]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[153:155]),
		.mem_out(sb_mux_size4_10_sram[0:2]),
		.mem_outb(sb_mux_size4_10_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_right_track_56 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[156:158]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[156:158]),
		.mem_out(sb_mux_size4_11_sram[0:2]),
		.mem_outb(sb_mux_size4_11_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_left_track_5 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[229:231]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[229:231]),
		.mem_out(sb_mux_size4_12_sram[0:2]),
		.mem_outb(sb_mux_size4_12_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_left_track_7 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[232:234]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[232:234]),
		.mem_out(sb_mux_size4_13_sram[0:2]),
		.mem_outb(sb_mux_size4_13_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_left_track_9 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[235:237]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[235:237]),
		.mem_out(sb_mux_size4_14_sram[0:2]),
		.mem_outb(sb_mux_size4_14_sram_inv[0:2]));

	sb_mux_size4_feedthrough_mem feedthrough_mem_left_track_11 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[238:240]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[238:240]),
		.mem_out(sb_mux_size4_15_sram[0:2]),
		.mem_outb(sb_mux_size4_15_sram_inv[0:2]));

	sb_mux_size3 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_a2f_o_0_, chanx_right_in[25], chanx_left_in[25]}),
		.sram(sb_mux_size3_0_sram[0:1]),
		.sram_inv(sb_mux_size3_0_sram_inv[0:1]),
		.out(chany_top_out[13]));

	sb_mux_size3 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_a2f_o_0_, chanx_right_in[26], chanx_left_in[26]}),
		.sram(sb_mux_size3_1_sram[0:1]),
		.sram_inv(sb_mux_size3_1_sram_inv[0:1]),
		.out(chany_top_out[14]));

	sb_mux_size3 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_a2f_o_0_, chanx_right_in[28], chanx_left_in[28]}),
		.sram(sb_mux_size3_2_sram[0:1]),
		.sram_inv(sb_mux_size3_2_sram_inv[0:1]),
		.out(chany_top_out[15]));

	sb_mux_size3 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_a2f_o_0_, chanx_right_in[29], chanx_left_in[29]}),
		.sram(sb_mux_size3_3_sram[0:1]),
		.sram_inv(sb_mux_size3_3_sram_inv[0:1]),
		.out(chany_top_out[16]));

	sb_mux_size3 mux_top_track_34 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_a2f_o_0_, chanx_right_in[30], chanx_left_in[30]}),
		.sram(sb_mux_size3_4_sram[0:1]),
		.sram_inv(sb_mux_size3_4_sram_inv[0:1]),
		.out(chany_top_out[17]));

	sb_mux_size3_feedthrough_mem feedthrough_mem_top_track_26 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[39:40]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[39:40]),
		.mem_out(sb_mux_size3_0_sram[0:1]),
		.mem_outb(sb_mux_size3_0_sram_inv[0:1]));

	sb_mux_size3_feedthrough_mem feedthrough_mem_top_track_28 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[41:42]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[41:42]),
		.mem_out(sb_mux_size3_1_sram[0:1]),
		.mem_outb(sb_mux_size3_1_sram_inv[0:1]));

	sb_mux_size3_feedthrough_mem feedthrough_mem_top_track_30 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[43:44]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[43:44]),
		.mem_out(sb_mux_size3_2_sram[0:1]),
		.mem_outb(sb_mux_size3_2_sram_inv[0:1]));

	sb_mux_size3_feedthrough_mem feedthrough_mem_top_track_32 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[45:46]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[45:46]),
		.mem_out(sb_mux_size3_3_sram[0:1]),
		.mem_outb(sb_mux_size3_3_sram_inv[0:1]));

	sb_mux_size3_feedthrough_mem feedthrough_mem_top_track_34 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[47:48]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[47:48]),
		.mem_out(sb_mux_size3_4_sram[0:1]),
		.mem_outb(sb_mux_size3_4_sram_inv[0:1]));

	sb_mux_size2 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_a2f_o_0_, chanx_left_in[31]}),
		.sram(sb_mux_size2_0_sram[0:1]),
		.sram_inv(sb_mux_size2_0_sram_inv[0:1]),
		.out(chany_top_out[19]));

	sb_mux_size2 mux_top_track_62 (
		.in({chanx_right_in[0], chanx_left_in[1]}),
		.sram(sb_mux_size2_1_sram[0:1]),
		.sram_inv(sb_mux_size2_1_sram_inv[0:1]),
		.out(chany_top_out[31]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_top_track_38 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[49:50]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[49:50]),
		.mem_out(sb_mux_size2_0_sram[0:1]),
		.mem_outb(sb_mux_size2_0_sram_inv[0:1]));

	sb_mux_size2_feedthrough_mem feedthrough_mem_top_track_62 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[51:52]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[51:52]),
		.mem_out(sb_mux_size2_1_sram[0:1]),
		.mem_outb(sb_mux_size2_1_sram_inv[0:1]));

	clk_mux_size3 mux_top_track_64 (
		.in({chanx_right_in[32], chany_bottom_in[0], chanx_left_in[32]}),
		.sram(clk_mux_size3_0_sram[0:1]),
		.sram_inv(clk_mux_size3_0_sram_inv[0:1]),
		.out(chany_top_out[32]));

	clk_mux_size3 mux_top_track_66 (
		.in({chanx_right_in[33], chany_bottom_in[1], chanx_left_in[33]}),
		.sram(clk_mux_size3_1_sram[0:1]),
		.sram_inv(clk_mux_size3_1_sram_inv[0:1]),
		.out(chany_top_out[33]));

	clk_mux_size3 mux_top_track_68 (
		.in({chanx_right_in[34], chany_bottom_in[2], chanx_left_in[34]}),
		.sram(clk_mux_size3_2_sram[0:1]),
		.sram_inv(clk_mux_size3_2_sram_inv[0:1]),
		.out(chany_top_out[34]));

	clk_mux_size3 mux_top_track_70 (
		.in({chanx_right_in[35], chany_bottom_in[3], chanx_left_in[35]}),
		.sram(clk_mux_size3_3_sram[0:1]),
		.sram_inv(clk_mux_size3_3_sram_inv[0:1]),
		.out(chany_top_out[35]));

	clk_mux_size3 mux_top_track_72 (
		.in({chanx_right_in[36], chany_bottom_in[4], chanx_left_in[36]}),
		.sram(clk_mux_size3_4_sram[0:1]),
		.sram_inv(clk_mux_size3_4_sram_inv[0:1]),
		.out(chany_top_out[36]));

	clk_mux_size3 mux_top_track_74 (
		.in({chanx_right_in[37], chany_bottom_in[5], chanx_left_in[37]}),
		.sram(clk_mux_size3_5_sram[0:1]),
		.sram_inv(clk_mux_size3_5_sram_inv[0:1]),
		.out(chany_top_out[37]));

	clk_mux_size3 mux_top_track_76 (
		.in({chanx_right_in[38], chany_bottom_in[6], chanx_left_in[38]}),
		.sram(clk_mux_size3_6_sram[0:1]),
		.sram_inv(clk_mux_size3_6_sram_inv[0:1]),
		.out(chany_top_out[38]));

	clk_mux_size3 mux_top_track_78 (
		.in({chanx_right_in[39], chany_bottom_in[7], chanx_left_in[39]}),
		.sram(clk_mux_size3_7_sram[0:1]),
		.sram_inv(clk_mux_size3_7_sram_inv[0:1]),
		.out(chany_top_out[39]));

	clk_mux_size3 mux_top_track_80 (
		.in({chanx_right_in[40], chany_bottom_in[8], chanx_left_in[40]}),
		.sram(clk_mux_size3_8_sram[0:1]),
		.sram_inv(clk_mux_size3_8_sram_inv[0:1]),
		.out(chany_top_out[40]));

	clk_mux_size3 mux_top_track_82 (
		.in({chanx_right_in[41], chany_bottom_in[9], chanx_left_in[41]}),
		.sram(clk_mux_size3_9_sram[0:1]),
		.sram_inv(clk_mux_size3_9_sram_inv[0:1]),
		.out(chany_top_out[41]));

	clk_mux_size3 mux_top_track_84 (
		.in({chanx_right_in[42], chany_bottom_in[10], chanx_left_in[42]}),
		.sram(clk_mux_size3_10_sram[0:1]),
		.sram_inv(clk_mux_size3_10_sram_inv[0:1]),
		.out(chany_top_out[42]));

	clk_mux_size3 mux_top_track_86 (
		.in({chanx_right_in[43], chany_bottom_in[11], chanx_left_in[43]}),
		.sram(clk_mux_size3_11_sram[0:1]),
		.sram_inv(clk_mux_size3_11_sram_inv[0:1]),
		.out(chany_top_out[43]));

	clk_mux_size3 mux_top_track_88 (
		.in({chanx_right_in[44], chany_bottom_in[12], chanx_left_in[44]}),
		.sram(clk_mux_size3_12_sram[0:1]),
		.sram_inv(clk_mux_size3_12_sram_inv[0:1]),
		.out(chany_top_out[44]));

	clk_mux_size3 mux_top_track_90 (
		.in({chanx_right_in[45], chany_bottom_in[13], chanx_left_in[45]}),
		.sram(clk_mux_size3_13_sram[0:1]),
		.sram_inv(clk_mux_size3_13_sram_inv[0:1]),
		.out(chany_top_out[45]));

	clk_mux_size3 mux_top_track_92 (
		.in({chanx_right_in[46], chany_bottom_in[14], chanx_left_in[46]}),
		.sram(clk_mux_size3_14_sram[0:1]),
		.sram_inv(clk_mux_size3_14_sram_inv[0:1]),
		.out(chany_top_out[46]));

	clk_mux_size3 mux_top_track_94 (
		.in({chanx_right_in[47], chany_bottom_in[15], chanx_left_in[47]}),
		.sram(clk_mux_size3_15_sram[0:1]),
		.sram_inv(clk_mux_size3_15_sram_inv[0:1]),
		.out(chany_top_out[47]));

	clk_mux_size3 mux_top_track_96 (
		.in({chanx_right_in[48], chany_bottom_in[16], chanx_left_in[48]}),
		.sram(clk_mux_size3_16_sram[0:1]),
		.sram_inv(clk_mux_size3_16_sram_inv[0:1]),
		.out(chany_top_out[48]));

	clk_mux_size3 mux_top_track_98 (
		.in({chanx_right_in[49], chany_bottom_in[17], chanx_left_in[49]}),
		.sram(clk_mux_size3_17_sram[0:1]),
		.sram_inv(clk_mux_size3_17_sram_inv[0:1]),
		.out(chany_top_out[49]));

	clk_mux_size3 mux_top_track_100 (
		.in({chanx_right_in[50], chany_bottom_in[18], chanx_left_in[50]}),
		.sram(clk_mux_size3_18_sram[0:1]),
		.sram_inv(clk_mux_size3_18_sram_inv[0:1]),
		.out(chany_top_out[50]));

	clk_mux_size3 mux_top_track_102 (
		.in({chanx_right_in[51], chany_bottom_in[19], chanx_left_in[51]}),
		.sram(clk_mux_size3_19_sram[0:1]),
		.sram_inv(clk_mux_size3_19_sram_inv[0:1]),
		.out(chany_top_out[51]));

	clk_mux_size3 mux_top_track_104 (
		.in({chanx_right_in[52], chany_bottom_in[20], chanx_left_in[52]}),
		.sram(clk_mux_size3_20_sram[0:1]),
		.sram_inv(clk_mux_size3_20_sram_inv[0:1]),
		.out(chany_top_out[52]));

	clk_mux_size3 mux_top_track_106 (
		.in({chanx_right_in[53], chany_bottom_in[21], chanx_left_in[53]}),
		.sram(clk_mux_size3_21_sram[0:1]),
		.sram_inv(clk_mux_size3_21_sram_inv[0:1]),
		.out(chany_top_out[53]));

	clk_mux_size3 mux_top_track_108 (
		.in({chanx_right_in[54], chany_bottom_in[22], chanx_left_in[54]}),
		.sram(clk_mux_size3_22_sram[0:1]),
		.sram_inv(clk_mux_size3_22_sram_inv[0:1]),
		.out(chany_top_out[54]));

	clk_mux_size3 mux_top_track_110 (
		.in({chanx_right_in[55], chany_bottom_in[23], chanx_left_in[55]}),
		.sram(clk_mux_size3_23_sram[0:1]),
		.sram_inv(clk_mux_size3_23_sram_inv[0:1]),
		.out(chany_top_out[55]));

	clk_mux_size3 mux_top_track_112 (
		.in({chanx_right_in[56], chany_bottom_in[24], chanx_left_in[56]}),
		.sram(clk_mux_size3_24_sram[0:1]),
		.sram_inv(clk_mux_size3_24_sram_inv[0:1]),
		.out(chany_top_out[56]));

	clk_mux_size3 mux_top_track_114 (
		.in({chanx_right_in[57], chany_bottom_in[25], chanx_left_in[57]}),
		.sram(clk_mux_size3_25_sram[0:1]),
		.sram_inv(clk_mux_size3_25_sram_inv[0:1]),
		.out(chany_top_out[57]));

	clk_mux_size3 mux_top_track_116 (
		.in({chanx_right_in[58], chany_bottom_in[26], chanx_left_in[58]}),
		.sram(clk_mux_size3_26_sram[0:1]),
		.sram_inv(clk_mux_size3_26_sram_inv[0:1]),
		.out(chany_top_out[58]));

	clk_mux_size3 mux_top_track_118 (
		.in({chanx_right_in[59], chany_bottom_in[27], chanx_left_in[59]}),
		.sram(clk_mux_size3_27_sram[0:1]),
		.sram_inv(clk_mux_size3_27_sram_inv[0:1]),
		.out(chany_top_out[59]));

	clk_mux_size3 mux_top_track_120 (
		.in({chanx_right_in[60], chany_bottom_in[28], chanx_left_in[60]}),
		.sram(clk_mux_size3_28_sram[0:1]),
		.sram_inv(clk_mux_size3_28_sram_inv[0:1]),
		.out(chany_top_out[60]));

	clk_mux_size3 mux_top_track_122 (
		.in({chanx_right_in[61], chany_bottom_in[29], chanx_left_in[61]}),
		.sram(clk_mux_size3_29_sram[0:1]),
		.sram_inv(clk_mux_size3_29_sram_inv[0:1]),
		.out(chany_top_out[61]));

	clk_mux_size3 mux_top_track_124 (
		.in({chanx_right_in[62], chany_bottom_in[30], chanx_left_in[62]}),
		.sram(clk_mux_size3_30_sram[0:1]),
		.sram_inv(clk_mux_size3_30_sram_inv[0:1]),
		.out(chany_top_out[62]));

	clk_mux_size3 mux_top_track_126 (
		.in({chanx_right_in[63], chany_bottom_in[31], chanx_left_in[63]}),
		.sram(clk_mux_size3_31_sram[0:1]),
		.sram_inv(clk_mux_size3_31_sram_inv[0:1]),
		.out(chany_top_out[63]));

	clk_mux_size3 mux_bottom_track_1 (
		.in({chany_top_in[32], chanx_right_in[32], chanx_left_in[32]}),
		.sram(clk_mux_size3_32_sram[0:1]),
		.sram_inv(clk_mux_size3_32_sram_inv[0:1]),
		.out(chany_bottom_out[0]));

	clk_mux_size3 mux_bottom_track_3 (
		.in({chany_top_in[33], chanx_right_in[33], chanx_left_in[33]}),
		.sram(clk_mux_size3_33_sram[0:1]),
		.sram_inv(clk_mux_size3_33_sram_inv[0:1]),
		.out(chany_bottom_out[1]));

	clk_mux_size3 mux_bottom_track_5 (
		.in({chany_top_in[34], chanx_right_in[34], chanx_left_in[34]}),
		.sram(clk_mux_size3_34_sram[0:1]),
		.sram_inv(clk_mux_size3_34_sram_inv[0:1]),
		.out(chany_bottom_out[2]));

	clk_mux_size3 mux_bottom_track_7 (
		.in({chany_top_in[35], chanx_right_in[35], chanx_left_in[35]}),
		.sram(clk_mux_size3_35_sram[0:1]),
		.sram_inv(clk_mux_size3_35_sram_inv[0:1]),
		.out(chany_bottom_out[3]));

	clk_mux_size3 mux_bottom_track_9 (
		.in({chany_top_in[36], chanx_right_in[36], chanx_left_in[36]}),
		.sram(clk_mux_size3_36_sram[0:1]),
		.sram_inv(clk_mux_size3_36_sram_inv[0:1]),
		.out(chany_bottom_out[4]));

	clk_mux_size3 mux_bottom_track_11 (
		.in({chany_top_in[37], chanx_right_in[37], chanx_left_in[37]}),
		.sram(clk_mux_size3_37_sram[0:1]),
		.sram_inv(clk_mux_size3_37_sram_inv[0:1]),
		.out(chany_bottom_out[5]));

	clk_mux_size3 mux_bottom_track_13 (
		.in({chany_top_in[38], chanx_right_in[38], chanx_left_in[38]}),
		.sram(clk_mux_size3_38_sram[0:1]),
		.sram_inv(clk_mux_size3_38_sram_inv[0:1]),
		.out(chany_bottom_out[6]));

	clk_mux_size3 mux_bottom_track_15 (
		.in({chany_top_in[39], chanx_right_in[39], chanx_left_in[39]}),
		.sram(clk_mux_size3_39_sram[0:1]),
		.sram_inv(clk_mux_size3_39_sram_inv[0:1]),
		.out(chany_bottom_out[7]));

	clk_mux_size3 mux_bottom_track_17 (
		.in({chany_top_in[40], chanx_right_in[40], chanx_left_in[40]}),
		.sram(clk_mux_size3_40_sram[0:1]),
		.sram_inv(clk_mux_size3_40_sram_inv[0:1]),
		.out(chany_bottom_out[8]));

	clk_mux_size3 mux_bottom_track_19 (
		.in({chany_top_in[41], chanx_right_in[41], chanx_left_in[41]}),
		.sram(clk_mux_size3_41_sram[0:1]),
		.sram_inv(clk_mux_size3_41_sram_inv[0:1]),
		.out(chany_bottom_out[9]));

	clk_mux_size3 mux_bottom_track_21 (
		.in({chany_top_in[42], chanx_right_in[42], chanx_left_in[42]}),
		.sram(clk_mux_size3_42_sram[0:1]),
		.sram_inv(clk_mux_size3_42_sram_inv[0:1]),
		.out(chany_bottom_out[10]));

	clk_mux_size3 mux_bottom_track_23 (
		.in({chany_top_in[43], chanx_right_in[43], chanx_left_in[43]}),
		.sram(clk_mux_size3_43_sram[0:1]),
		.sram_inv(clk_mux_size3_43_sram_inv[0:1]),
		.out(chany_bottom_out[11]));

	clk_mux_size3 mux_bottom_track_25 (
		.in({chany_top_in[44], chanx_right_in[44], chanx_left_in[44]}),
		.sram(clk_mux_size3_44_sram[0:1]),
		.sram_inv(clk_mux_size3_44_sram_inv[0:1]),
		.out(chany_bottom_out[12]));

	clk_mux_size3 mux_bottom_track_27 (
		.in({chany_top_in[45], chanx_right_in[45], chanx_left_in[45]}),
		.sram(clk_mux_size3_45_sram[0:1]),
		.sram_inv(clk_mux_size3_45_sram_inv[0:1]),
		.out(chany_bottom_out[13]));

	clk_mux_size3 mux_bottom_track_29 (
		.in({chany_top_in[46], chanx_right_in[46], chanx_left_in[46]}),
		.sram(clk_mux_size3_46_sram[0:1]),
		.sram_inv(clk_mux_size3_46_sram_inv[0:1]),
		.out(chany_bottom_out[14]));

	clk_mux_size3 mux_bottom_track_31 (
		.in({chany_top_in[47], chanx_right_in[47], chanx_left_in[47]}),
		.sram(clk_mux_size3_47_sram[0:1]),
		.sram_inv(clk_mux_size3_47_sram_inv[0:1]),
		.out(chany_bottom_out[15]));

	clk_mux_size3 mux_bottom_track_33 (
		.in({chany_top_in[48], chanx_right_in[48], chanx_left_in[48]}),
		.sram(clk_mux_size3_48_sram[0:1]),
		.sram_inv(clk_mux_size3_48_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	clk_mux_size3 mux_bottom_track_35 (
		.in({chany_top_in[49], chanx_right_in[49], chanx_left_in[49]}),
		.sram(clk_mux_size3_49_sram[0:1]),
		.sram_inv(clk_mux_size3_49_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	clk_mux_size3 mux_bottom_track_37 (
		.in({chany_top_in[50], chanx_right_in[50], chanx_left_in[50]}),
		.sram(clk_mux_size3_50_sram[0:1]),
		.sram_inv(clk_mux_size3_50_sram_inv[0:1]),
		.out(chany_bottom_out[18]));

	clk_mux_size3 mux_bottom_track_39 (
		.in({chany_top_in[51], chanx_right_in[51], chanx_left_in[51]}),
		.sram(clk_mux_size3_51_sram[0:1]),
		.sram_inv(clk_mux_size3_51_sram_inv[0:1]),
		.out(chany_bottom_out[19]));

	clk_mux_size3 mux_bottom_track_41 (
		.in({chany_top_in[52], chanx_right_in[52], chanx_left_in[52]}),
		.sram(clk_mux_size3_52_sram[0:1]),
		.sram_inv(clk_mux_size3_52_sram_inv[0:1]),
		.out(chany_bottom_out[20]));

	clk_mux_size3 mux_bottom_track_43 (
		.in({chany_top_in[53], chanx_right_in[53], chanx_left_in[53]}),
		.sram(clk_mux_size3_53_sram[0:1]),
		.sram_inv(clk_mux_size3_53_sram_inv[0:1]),
		.out(chany_bottom_out[21]));

	clk_mux_size3 mux_bottom_track_45 (
		.in({chany_top_in[54], chanx_right_in[54], chanx_left_in[54]}),
		.sram(clk_mux_size3_54_sram[0:1]),
		.sram_inv(clk_mux_size3_54_sram_inv[0:1]),
		.out(chany_bottom_out[22]));

	clk_mux_size3 mux_bottom_track_47 (
		.in({chany_top_in[55], chanx_right_in[55], chanx_left_in[55]}),
		.sram(clk_mux_size3_55_sram[0:1]),
		.sram_inv(clk_mux_size3_55_sram_inv[0:1]),
		.out(chany_bottom_out[23]));

	clk_mux_size3 mux_bottom_track_49 (
		.in({chany_top_in[56], chanx_right_in[56], chanx_left_in[56]}),
		.sram(clk_mux_size3_56_sram[0:1]),
		.sram_inv(clk_mux_size3_56_sram_inv[0:1]),
		.out(chany_bottom_out[24]));

	clk_mux_size3 mux_bottom_track_51 (
		.in({chany_top_in[57], chanx_right_in[57], chanx_left_in[57]}),
		.sram(clk_mux_size3_57_sram[0:1]),
		.sram_inv(clk_mux_size3_57_sram_inv[0:1]),
		.out(chany_bottom_out[25]));

	clk_mux_size3 mux_bottom_track_53 (
		.in({chany_top_in[58], chanx_right_in[58], chanx_left_in[58]}),
		.sram(clk_mux_size3_58_sram[0:1]),
		.sram_inv(clk_mux_size3_58_sram_inv[0:1]),
		.out(chany_bottom_out[26]));

	clk_mux_size3 mux_bottom_track_55 (
		.in({chany_top_in[59], chanx_right_in[59], chanx_left_in[59]}),
		.sram(clk_mux_size3_59_sram[0:1]),
		.sram_inv(clk_mux_size3_59_sram_inv[0:1]),
		.out(chany_bottom_out[27]));

	clk_mux_size3 mux_bottom_track_57 (
		.in({chany_top_in[60], chanx_right_in[60], chanx_left_in[60]}),
		.sram(clk_mux_size3_60_sram[0:1]),
		.sram_inv(clk_mux_size3_60_sram_inv[0:1]),
		.out(chany_bottom_out[28]));

	clk_mux_size3 mux_bottom_track_59 (
		.in({chany_top_in[61], chanx_right_in[61], chanx_left_in[61]}),
		.sram(clk_mux_size3_61_sram[0:1]),
		.sram_inv(clk_mux_size3_61_sram_inv[0:1]),
		.out(chany_bottom_out[29]));

	clk_mux_size3 mux_bottom_track_61 (
		.in({chany_top_in[62], chanx_right_in[62], chanx_left_in[62]}),
		.sram(clk_mux_size3_62_sram[0:1]),
		.sram_inv(clk_mux_size3_62_sram_inv[0:1]),
		.out(chany_bottom_out[30]));

	clk_mux_size3 mux_bottom_track_63 (
		.in({chany_top_in[63], chanx_right_in[63], chanx_left_in[63]}),
		.sram(clk_mux_size3_63_sram[0:1]),
		.sram_inv(clk_mux_size3_63_sram_inv[0:1]),
		.out(chany_bottom_out[31]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_64 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[53:54]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[53:54]),
		.mem_out(clk_mux_size3_0_sram[0:1]),
		.mem_outb(clk_mux_size3_0_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_66 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[55:56]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[55:56]),
		.mem_out(clk_mux_size3_1_sram[0:1]),
		.mem_outb(clk_mux_size3_1_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_68 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[57:58]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[57:58]),
		.mem_out(clk_mux_size3_2_sram[0:1]),
		.mem_outb(clk_mux_size3_2_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_70 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[59:60]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[59:60]),
		.mem_out(clk_mux_size3_3_sram[0:1]),
		.mem_outb(clk_mux_size3_3_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_72 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[61:62]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[61:62]),
		.mem_out(clk_mux_size3_4_sram[0:1]),
		.mem_outb(clk_mux_size3_4_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_74 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[63:64]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[63:64]),
		.mem_out(clk_mux_size3_5_sram[0:1]),
		.mem_outb(clk_mux_size3_5_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_76 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[65:66]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[65:66]),
		.mem_out(clk_mux_size3_6_sram[0:1]),
		.mem_outb(clk_mux_size3_6_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_78 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[67:68]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[67:68]),
		.mem_out(clk_mux_size3_7_sram[0:1]),
		.mem_outb(clk_mux_size3_7_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_80 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[69:70]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[69:70]),
		.mem_out(clk_mux_size3_8_sram[0:1]),
		.mem_outb(clk_mux_size3_8_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_82 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[71:72]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[71:72]),
		.mem_out(clk_mux_size3_9_sram[0:1]),
		.mem_outb(clk_mux_size3_9_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_84 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[73:74]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[73:74]),
		.mem_out(clk_mux_size3_10_sram[0:1]),
		.mem_outb(clk_mux_size3_10_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_86 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[75:76]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[75:76]),
		.mem_out(clk_mux_size3_11_sram[0:1]),
		.mem_outb(clk_mux_size3_11_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_88 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[77:78]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[77:78]),
		.mem_out(clk_mux_size3_12_sram[0:1]),
		.mem_outb(clk_mux_size3_12_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_90 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[79:80]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[79:80]),
		.mem_out(clk_mux_size3_13_sram[0:1]),
		.mem_outb(clk_mux_size3_13_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_92 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[81:82]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[81:82]),
		.mem_out(clk_mux_size3_14_sram[0:1]),
		.mem_outb(clk_mux_size3_14_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_94 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[83:84]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[83:84]),
		.mem_out(clk_mux_size3_15_sram[0:1]),
		.mem_outb(clk_mux_size3_15_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_96 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[85:86]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[85:86]),
		.mem_out(clk_mux_size3_16_sram[0:1]),
		.mem_outb(clk_mux_size3_16_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_98 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[87:88]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[87:88]),
		.mem_out(clk_mux_size3_17_sram[0:1]),
		.mem_outb(clk_mux_size3_17_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_100 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[89:90]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[89:90]),
		.mem_out(clk_mux_size3_18_sram[0:1]),
		.mem_outb(clk_mux_size3_18_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_102 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[91:92]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[91:92]),
		.mem_out(clk_mux_size3_19_sram[0:1]),
		.mem_outb(clk_mux_size3_19_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_104 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[93:94]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[93:94]),
		.mem_out(clk_mux_size3_20_sram[0:1]),
		.mem_outb(clk_mux_size3_20_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_106 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[95:96]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[95:96]),
		.mem_out(clk_mux_size3_21_sram[0:1]),
		.mem_outb(clk_mux_size3_21_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_108 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[97:98]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[97:98]),
		.mem_out(clk_mux_size3_22_sram[0:1]),
		.mem_outb(clk_mux_size3_22_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_110 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[99:100]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[99:100]),
		.mem_out(clk_mux_size3_23_sram[0:1]),
		.mem_outb(clk_mux_size3_23_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_112 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[101:102]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[101:102]),
		.mem_out(clk_mux_size3_24_sram[0:1]),
		.mem_outb(clk_mux_size3_24_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_114 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[103:104]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[103:104]),
		.mem_out(clk_mux_size3_25_sram[0:1]),
		.mem_outb(clk_mux_size3_25_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_116 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[105:106]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[105:106]),
		.mem_out(clk_mux_size3_26_sram[0:1]),
		.mem_outb(clk_mux_size3_26_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_118 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[107:108]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[107:108]),
		.mem_out(clk_mux_size3_27_sram[0:1]),
		.mem_outb(clk_mux_size3_27_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_120 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[109:110]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[109:110]),
		.mem_out(clk_mux_size3_28_sram[0:1]),
		.mem_outb(clk_mux_size3_28_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_122 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[111:112]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[111:112]),
		.mem_out(clk_mux_size3_29_sram[0:1]),
		.mem_outb(clk_mux_size3_29_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_124 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[113:114]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[113:114]),
		.mem_out(clk_mux_size3_30_sram[0:1]),
		.mem_outb(clk_mux_size3_30_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_top_track_126 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[115:116]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[115:116]),
		.mem_out(clk_mux_size3_31_sram[0:1]),
		.mem_outb(clk_mux_size3_31_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_1 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[159:160]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[159:160]),
		.mem_out(clk_mux_size3_32_sram[0:1]),
		.mem_outb(clk_mux_size3_32_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_3 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[161:162]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[161:162]),
		.mem_out(clk_mux_size3_33_sram[0:1]),
		.mem_outb(clk_mux_size3_33_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_5 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[163:164]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[163:164]),
		.mem_out(clk_mux_size3_34_sram[0:1]),
		.mem_outb(clk_mux_size3_34_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_7 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[165:166]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[165:166]),
		.mem_out(clk_mux_size3_35_sram[0:1]),
		.mem_outb(clk_mux_size3_35_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_9 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[167:168]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[167:168]),
		.mem_out(clk_mux_size3_36_sram[0:1]),
		.mem_outb(clk_mux_size3_36_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_11 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[169:170]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[169:170]),
		.mem_out(clk_mux_size3_37_sram[0:1]),
		.mem_outb(clk_mux_size3_37_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_13 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[171:172]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[171:172]),
		.mem_out(clk_mux_size3_38_sram[0:1]),
		.mem_outb(clk_mux_size3_38_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_15 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[173:174]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[173:174]),
		.mem_out(clk_mux_size3_39_sram[0:1]),
		.mem_outb(clk_mux_size3_39_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_17 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[175:176]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[175:176]),
		.mem_out(clk_mux_size3_40_sram[0:1]),
		.mem_outb(clk_mux_size3_40_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_19 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[177:178]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[177:178]),
		.mem_out(clk_mux_size3_41_sram[0:1]),
		.mem_outb(clk_mux_size3_41_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_21 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[179:180]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[179:180]),
		.mem_out(clk_mux_size3_42_sram[0:1]),
		.mem_outb(clk_mux_size3_42_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_23 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[181:182]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[181:182]),
		.mem_out(clk_mux_size3_43_sram[0:1]),
		.mem_outb(clk_mux_size3_43_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_25 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[183:184]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[183:184]),
		.mem_out(clk_mux_size3_44_sram[0:1]),
		.mem_outb(clk_mux_size3_44_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_27 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[185:186]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[185:186]),
		.mem_out(clk_mux_size3_45_sram[0:1]),
		.mem_outb(clk_mux_size3_45_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_29 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[187:188]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[187:188]),
		.mem_out(clk_mux_size3_46_sram[0:1]),
		.mem_outb(clk_mux_size3_46_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_31 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[189:190]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[189:190]),
		.mem_out(clk_mux_size3_47_sram[0:1]),
		.mem_outb(clk_mux_size3_47_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_33 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[191:192]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[191:192]),
		.mem_out(clk_mux_size3_48_sram[0:1]),
		.mem_outb(clk_mux_size3_48_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_35 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[193:194]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[193:194]),
		.mem_out(clk_mux_size3_49_sram[0:1]),
		.mem_outb(clk_mux_size3_49_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_37 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[195:196]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[195:196]),
		.mem_out(clk_mux_size3_50_sram[0:1]),
		.mem_outb(clk_mux_size3_50_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_39 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[197:198]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[197:198]),
		.mem_out(clk_mux_size3_51_sram[0:1]),
		.mem_outb(clk_mux_size3_51_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_41 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[199:200]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[199:200]),
		.mem_out(clk_mux_size3_52_sram[0:1]),
		.mem_outb(clk_mux_size3_52_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_43 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[201:202]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[201:202]),
		.mem_out(clk_mux_size3_53_sram[0:1]),
		.mem_outb(clk_mux_size3_53_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_45 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[203:204]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[203:204]),
		.mem_out(clk_mux_size3_54_sram[0:1]),
		.mem_outb(clk_mux_size3_54_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_47 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[205:206]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[205:206]),
		.mem_out(clk_mux_size3_55_sram[0:1]),
		.mem_outb(clk_mux_size3_55_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_49 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[207:208]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[207:208]),
		.mem_out(clk_mux_size3_56_sram[0:1]),
		.mem_outb(clk_mux_size3_56_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_51 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[209:210]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[209:210]),
		.mem_out(clk_mux_size3_57_sram[0:1]),
		.mem_outb(clk_mux_size3_57_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_53 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[211:212]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[211:212]),
		.mem_out(clk_mux_size3_58_sram[0:1]),
		.mem_outb(clk_mux_size3_58_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_55 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[213:214]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[213:214]),
		.mem_out(clk_mux_size3_59_sram[0:1]),
		.mem_outb(clk_mux_size3_59_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_57 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[215:216]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[215:216]),
		.mem_out(clk_mux_size3_60_sram[0:1]),
		.mem_outb(clk_mux_size3_60_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_59 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[217:218]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[217:218]),
		.mem_out(clk_mux_size3_61_sram[0:1]),
		.mem_outb(clk_mux_size3_61_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_61 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[219:220]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[219:220]),
		.mem_out(clk_mux_size3_62_sram[0:1]),
		.mem_outb(clk_mux_size3_62_sram_inv[0:1]));

	clk_mux_size3_feedthrough_mem feedthrough_mem_bottom_track_63 (
		.feedthrough_mem_in(sb_0__config_group_mem_size265_0_mem_out[221:222]),
		.feedthrough_mem_inb(sb_0__config_group_mem_size265_0_mem_outb[221:222]),
		.mem_out(clk_mux_size3_63_sram[0:1]),
		.mem_outb(clk_mux_size3_63_sram_inv[0:1]));

	sb_0__config_group_mem_size265 sb_0__config_group_mem_size265 (
		.config_enable(config_enable),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.mem_out(sb_0__config_group_mem_size265_0_mem_out[0:264]),
		.mem_outb(sb_0__config_group_mem_size265_0_mem_outb[0:264]),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for sb_0_ -----



